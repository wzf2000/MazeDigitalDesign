module intersection
#parameter( wall = 0)
(
    input wire clk,
    input wire signed [9:0] dir,    // * 2 ^ 8
    input wire signed [9:0] ori,    // * 2 ^ 0
    output reg signed [18:0] p      // * 2 ^ 0
);

localparam [0:511][8:0] inverse = {
    9'b111111111,
    9'b111111111,
    9'd100000000,
    9'd010101011,
    9'd010000000,
    9'd001100110,
    9'd001010101,
    9'd001001001,
    9'd001000000,
    9'd000111001,
    9'd000110011,
    9'd000101111,
    9'd000101011,
    9'd000100111,
    9'd000100101,
    9'd000100010,
    9'd000100000,
    9'd000011110,
    9'd000011100,
    9'd000011011,
    9'd000011010,
    9'd000011000,
    9'd000010111,
    9'd000010110,
    9'd000010101,
    9'd000010100,
    9'd000010100,
    9'd000010011,
    9'd000010010,
    9'd000010010,
    9'd000010001,
    9'd000010001,
    9'd000010000,
    9'd000010000,
    9'd000001111,
    9'd000001111,
    9'd000001110,
    9'd000001110,
    9'd000001101,
    9'd000001101,
    9'd000001101,
    9'd000001100,
    9'd000001100,
    9'd000001100,
    9'd000001100,
    9'd000001011,
    9'd000001011,
    9'd000001011,
    9'd000001011,
    9'd000001010,
    9'd000001010,
    9'd000001010,
    9'd000001010,
    9'd000001010,
    9'd000001001,
    9'd000001001,
    9'd000001001,
    9'd000001001,
    9'd000001001,
    9'd000001001,
    9'd000001001,
    9'd000001000,
    9'd000001000,
    9'd000001000,
    9'd000001000,
    9'd000001000,
    9'd000001000,
    9'd000001000,
    9'd000001000,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000111,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000110,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000101,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000100,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000011,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000010,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001,
    9'd000000001
};

wire less;
wire sign;

assign less = (wall << 6) < ori;
assign sign = dir[9] ^ less;

always @(posedge clk) begin
    if (dir[8:0] == 10'd0) begin
        p <= 19'b1111111111111111111;
    end
    else begin
        if (sign)
            p <= 19'b1111111111111111111;
        else begin
            p[18] <= 1'b0;
            p[17:0] <= ((less ? (ori - (wall << 6)) : ((wall << 6) - ori)) * inverse[dir[8:0]]) >> 1;
        end
    end
end

endmodule
