module intersection
#(parameter wall = 0)
(
    input wire clk,
    input wire signed [9:0] dir,    // * 2 ^ 8
    input wire signed [9:0] ori,    // * 2 ^ 0
    output reg signed [18:0] p      // * 2 ^ 0
);

localparam [0:511][15:0] inverse = {
	16'b1111111111111111,
	16'b1111111111111111,
	16'b1000000000000000,
	16'b0101010101010101,
	16'b0100000000000000,
	16'b0011001100110011,
	16'b0010101010101011,
	16'b0010010010010010,
	16'b0010000000000000,
	16'b0001110001110010,
	16'b0001100110011010,
	16'b0001011101000110,
	16'b0001010101010101,
	16'b0001001110110001,
	16'b0001001001001001,
	16'b0001000100010001,
	16'b0001000000000000,
	16'b0000111100001111,
	16'b0000111000111001,
	16'b0000110101111001,
	16'b0000110011001101,
	16'b0000110000110001,
	16'b0000101110100011,
	16'b0000101100100001,
	16'b0000101010101011,
	16'b0000101000111101,
	16'b0000100111011001,
	16'b0000100101111011,
	16'b0000100100100101,
	16'b0000100011010100,
	16'b0000100010001001,
	16'b0000100001000010,
	16'b0000100000000000,
	16'b0000011111000010,
	16'b0000011110001000,
	16'b0000011101010000,
	16'b0000011100011100,
	16'b0000011011101011,
	16'b0000011010111101,
	16'b0000011010010000,
	16'b0000011001100110,
	16'b0000011000111110,
	16'b0000011000011000,
	16'b0000010111110100,
	16'b0000010111010001,
	16'b0000010110110000,
	16'b0000010110010001,
	16'b0000010101110010,
	16'b0000010101010101,
	16'b0000010100111001,
	16'b0000010100011111,
	16'b0000010100000101,
	16'b0000010011101100,
	16'b0000010011010101,
	16'b0000010010111110,
	16'b0000010010101000,
	16'b0000010010010010,
	16'b0000010001111110,
	16'b0000010001101010,
	16'b0000010001010111,
	16'b0000010001000100,
	16'b0000010000110010,
	16'b0000010000100001,
	16'b0000010000010000,
	16'b0000010000000000,
	16'b0000001111110000,
	16'b0000001111100001,
	16'b0000001111010010,
	16'b0000001111000100,
	16'b0000001110110110,
	16'b0000001110101000,
	16'b0000001110011011,
	16'b0000001110001110,
	16'b0000001110000010,
	16'b0000001101110110,
	16'b0000001101101010,
	16'b0000001101011110,
	16'b0000001101010011,
	16'b0000001101001000,
	16'b0000001100111110,
	16'b0000001100110011,
	16'b0000001100101001,
	16'b0000001100011111,
	16'b0000001100010110,
	16'b0000001100001100,
	16'b0000001100000011,
	16'b0000001011111010,
	16'b0000001011110001,
	16'b0000001011101001,
	16'b0000001011100000,
	16'b0000001011011000,
	16'b0000001011010000,
	16'b0000001011001000,
	16'b0000001011000001,
	16'b0000001010111001,
	16'b0000001010110010,
	16'b0000001010101011,
	16'b0000001010100100,
	16'b0000001010011101,
	16'b0000001010010110,
	16'b0000001010001111,
	16'b0000001010001001,
	16'b0000001010000011,
	16'b0000001001111100,
	16'b0000001001110110,
	16'b0000001001110000,
	16'b0000001001101010,
	16'b0000001001100100,
	16'b0000001001011111,
	16'b0000001001011001,
	16'b0000001001010100,
	16'b0000001001001110,
	16'b0000001001001001,
	16'b0000001001000100,
	16'b0000001000111111,
	16'b0000001000111010,
	16'b0000001000110101,
	16'b0000001000110000,
	16'b0000001000101011,
	16'b0000001000100111,
	16'b0000001000100010,
	16'b0000001000011110,
	16'b0000001000011001,
	16'b0000001000010101,
	16'b0000001000010001,
	16'b0000001000001100,
	16'b0000001000001000,
	16'b0000001000000100,
	16'b0000001000000000,
	16'b0000000111111100,
	16'b0000000111111000,
	16'b0000000111110100,
	16'b0000000111110000,
	16'b0000000111101101,
	16'b0000000111101001,
	16'b0000000111100101,
	16'b0000000111100010,
	16'b0000000111011110,
	16'b0000000111011011,
	16'b0000000111010111,
	16'b0000000111010100,
	16'b0000000111010001,
	16'b0000000111001110,
	16'b0000000111001010,
	16'b0000000111000111,
	16'b0000000111000100,
	16'b0000000111000001,
	16'b0000000110111110,
	16'b0000000110111011,
	16'b0000000110111000,
	16'b0000000110110101,
	16'b0000000110110010,
	16'b0000000110101111,
	16'b0000000110101100,
	16'b0000000110101010,
	16'b0000000110100111,
	16'b0000000110100100,
	16'b0000000110100001,
	16'b0000000110011111,
	16'b0000000110011100,
	16'b0000000110011010,
	16'b0000000110010111,
	16'b0000000110010101,
	16'b0000000110010010,
	16'b0000000110010000,
	16'b0000000110001101,
	16'b0000000110001011,
	16'b0000000110001000,
	16'b0000000110000110,
	16'b0000000110000100,
	16'b0000000110000010,
	16'b0000000101111111,
	16'b0000000101111101,
	16'b0000000101111011,
	16'b0000000101111001,
	16'b0000000101110110,
	16'b0000000101110100,
	16'b0000000101110010,
	16'b0000000101110000,
	16'b0000000101101110,
	16'b0000000101101100,
	16'b0000000101101010,
	16'b0000000101101000,
	16'b0000000101100110,
	16'b0000000101100100,
	16'b0000000101100010,
	16'b0000000101100000,
	16'b0000000101011110,
	16'b0000000101011101,
	16'b0000000101011011,
	16'b0000000101011001,
	16'b0000000101010111,
	16'b0000000101010101,
	16'b0000000101010100,
	16'b0000000101010010,
	16'b0000000101010000,
	16'b0000000101001110,
	16'b0000000101001101,
	16'b0000000101001011,
	16'b0000000101001001,
	16'b0000000101001000,
	16'b0000000101000110,
	16'b0000000101000100,
	16'b0000000101000011,
	16'b0000000101000001,
	16'b0000000101000000,
	16'b0000000100111110,
	16'b0000000100111101,
	16'b0000000100111011,
	16'b0000000100111010,
	16'b0000000100111000,
	16'b0000000100110111,
	16'b0000000100110101,
	16'b0000000100110100,
	16'b0000000100110010,
	16'b0000000100110001,
	16'b0000000100101111,
	16'b0000000100101110,
	16'b0000000100101101,
	16'b0000000100101011,
	16'b0000000100101010,
	16'b0000000100101001,
	16'b0000000100100111,
	16'b0000000100100110,
	16'b0000000100100101,
	16'b0000000100100011,
	16'b0000000100100010,
	16'b0000000100100001,
	16'b0000000100011111,
	16'b0000000100011110,
	16'b0000000100011101,
	16'b0000000100011100,
	16'b0000000100011010,
	16'b0000000100011001,
	16'b0000000100011000,
	16'b0000000100010111,
	16'b0000000100010110,
	16'b0000000100010101,
	16'b0000000100010011,
	16'b0000000100010010,
	16'b0000000100010001,
	16'b0000000100010000,
	16'b0000000100001111,
	16'b0000000100001110,
	16'b0000000100001101,
	16'b0000000100001011,
	16'b0000000100001010,
	16'b0000000100001001,
	16'b0000000100001000,
	16'b0000000100000111,
	16'b0000000100000110,
	16'b0000000100000101,
	16'b0000000100000100,
	16'b0000000100000011,
	16'b0000000100000010,
	16'b0000000100000001,
	16'b0000000100000000,
	16'b0000000011111111,
	16'b0000000011111110,
	16'b0000000011111101,
	16'b0000000011111100,
	16'b0000000011111011,
	16'b0000000011111010,
	16'b0000000011111001,
	16'b0000000011111000,
	16'b0000000011110111,
	16'b0000000011110110,
	16'b0000000011110101,
	16'b0000000011110101,
	16'b0000000011110100,
	16'b0000000011110011,
	16'b0000000011110010,
	16'b0000000011110001,
	16'b0000000011110000,
	16'b0000000011101111,
	16'b0000000011101110,
	16'b0000000011101101,
	16'b0000000011101101,
	16'b0000000011101100,
	16'b0000000011101011,
	16'b0000000011101010,
	16'b0000000011101001,
	16'b0000000011101000,
	16'b0000000011101000,
	16'b0000000011100111,
	16'b0000000011100110,
	16'b0000000011100101,
	16'b0000000011100100,
	16'b0000000011100100,
	16'b0000000011100011,
	16'b0000000011100010,
	16'b0000000011100001,
	16'b0000000011100000,
	16'b0000000011100000,
	16'b0000000011011111,
	16'b0000000011011110,
	16'b0000000011011101,
	16'b0000000011011101,
	16'b0000000011011100,
	16'b0000000011011011,
	16'b0000000011011010,
	16'b0000000011011010,
	16'b0000000011011001,
	16'b0000000011011000,
	16'b0000000011011000,
	16'b0000000011010111,
	16'b0000000011010110,
	16'b0000000011010101,
	16'b0000000011010101,
	16'b0000000011010100,
	16'b0000000011010011,
	16'b0000000011010011,
	16'b0000000011010010,
	16'b0000000011010001,
	16'b0000000011010001,
	16'b0000000011010000,
	16'b0000000011001111,
	16'b0000000011001111,
	16'b0000000011001110,
	16'b0000000011001101,
	16'b0000000011001101,
	16'b0000000011001100,
	16'b0000000011001100,
	16'b0000000011001011,
	16'b0000000011001010,
	16'b0000000011001010,
	16'b0000000011001001,
	16'b0000000011001000,
	16'b0000000011001000,
	16'b0000000011000111,
	16'b0000000011000111,
	16'b0000000011000110,
	16'b0000000011000101,
	16'b0000000011000101,
	16'b0000000011000100,
	16'b0000000011000100,
	16'b0000000011000011,
	16'b0000000011000010,
	16'b0000000011000010,
	16'b0000000011000001,
	16'b0000000011000001,
	16'b0000000011000000,
	16'b0000000011000000,
	16'b0000000010111111,
	16'b0000000010111111,
	16'b0000000010111110,
	16'b0000000010111101,
	16'b0000000010111101,
	16'b0000000010111100,
	16'b0000000010111100,
	16'b0000000010111011,
	16'b0000000010111011,
	16'b0000000010111010,
	16'b0000000010111010,
	16'b0000000010111001,
	16'b0000000010111001,
	16'b0000000010111000,
	16'b0000000010111000,
	16'b0000000010110111,
	16'b0000000010110111,
	16'b0000000010110110,
	16'b0000000010110110,
	16'b0000000010110101,
	16'b0000000010110101,
	16'b0000000010110100,
	16'b0000000010110100,
	16'b0000000010110011,
	16'b0000000010110011,
	16'b0000000010110010,
	16'b0000000010110010,
	16'b0000000010110001,
	16'b0000000010110001,
	16'b0000000010110000,
	16'b0000000010110000,
	16'b0000000010101111,
	16'b0000000010101111,
	16'b0000000010101110,
	16'b0000000010101110,
	16'b0000000010101101,
	16'b0000000010101101,
	16'b0000000010101100,
	16'b0000000010101100,
	16'b0000000010101100,
	16'b0000000010101011,
	16'b0000000010101011,
	16'b0000000010101010,
	16'b0000000010101010,
	16'b0000000010101001,
	16'b0000000010101001,
	16'b0000000010101000,
	16'b0000000010101000,
	16'b0000000010101000,
	16'b0000000010100111,
	16'b0000000010100111,
	16'b0000000010100110,
	16'b0000000010100110,
	16'b0000000010100101,
	16'b0000000010100101,
	16'b0000000010100101,
	16'b0000000010100100,
	16'b0000000010100100,
	16'b0000000010100011,
	16'b0000000010100011,
	16'b0000000010100011,
	16'b0000000010100010,
	16'b0000000010100010,
	16'b0000000010100001,
	16'b0000000010100001,
	16'b0000000010100001,
	16'b0000000010100000,
	16'b0000000010100000,
	16'b0000000010011111,
	16'b0000000010011111,
	16'b0000000010011111,
	16'b0000000010011110,
	16'b0000000010011110,
	16'b0000000010011110,
	16'b0000000010011101,
	16'b0000000010011101,
	16'b0000000010011100,
	16'b0000000010011100,
	16'b0000000010011100,
	16'b0000000010011011,
	16'b0000000010011011,
	16'b0000000010011011,
	16'b0000000010011010,
	16'b0000000010011010,
	16'b0000000010011001,
	16'b0000000010011001,
	16'b0000000010011001,
	16'b0000000010011000,
	16'b0000000010011000,
	16'b0000000010011000,
	16'b0000000010010111,
	16'b0000000010010111,
	16'b0000000010010111,
	16'b0000000010010110,
	16'b0000000010010110,
	16'b0000000010010110,
	16'b0000000010010101,
	16'b0000000010010101,
	16'b0000000010010101,
	16'b0000000010010100,
	16'b0000000010010100,
	16'b0000000010010100,
	16'b0000000010010011,
	16'b0000000010010011,
	16'b0000000010010011,
	16'b0000000010010010,
	16'b0000000010010010,
	16'b0000000010010010,
	16'b0000000010010001,
	16'b0000000010010001,
	16'b0000000010010001,
	16'b0000000010010000,
	16'b0000000010010000,
	16'b0000000010010000,
	16'b0000000010001111,
	16'b0000000010001111,
	16'b0000000010001111,
	16'b0000000010001110,
	16'b0000000010001110,
	16'b0000000010001110,
	16'b0000000010001110,
	16'b0000000010001101,
	16'b0000000010001101,
	16'b0000000010001101,
	16'b0000000010001100,
	16'b0000000010001100,
	16'b0000000010001100,
	16'b0000000010001011,
	16'b0000000010001011,
	16'b0000000010001011,
	16'b0000000010001011,
	16'b0000000010001010,
	16'b0000000010001010,
	16'b0000000010001010,
	16'b0000000010001001,
	16'b0000000010001001,
	16'b0000000010001001,
	16'b0000000010001001,
	16'b0000000010001000,
	16'b0000000010001000,
	16'b0000000010001000,
	16'b0000000010000111,
	16'b0000000010000111,
	16'b0000000010000111,
	16'b0000000010000111,
	16'b0000000010000110,
	16'b0000000010000110,
	16'b0000000010000110,
	16'b0000000010000101,
	16'b0000000010000101,
	16'b0000000010000101,
	16'b0000000010000101,
	16'b0000000010000100,
	16'b0000000010000100,
	16'b0000000010000100,
	16'b0000000010000100,
	16'b0000000010000011,
	16'b0000000010000011,
	16'b0000000010000011,
	16'b0000000010000011,
	16'b0000000010000010,
	16'b0000000010000010,
	16'b0000000010000010,
	16'b0000000010000010,
	16'b0000000010000001,
	16'b0000000010000001,
	16'b0000000010000001,
	16'b0000000010000001,
	16'b0000000010000000
};

wire less;
wire sign;
wire signed [9:0] abs_dir;

assign less = (wall << 6) < ori;
assign sign = dir[9] ^ less;
assign abs_dir = dir[9] ? -dir : dir;

always @(posedge clk) begin
    if (dir[8:0] == 10'd0) begin
        p <= 19'b1111111111111111111;
    end
    else begin
        if (sign)
            p <= 19'b1111111111111111111;
        else begin
            p[18] <= 1'b0;
            p[17:0] <= ((less ? (ori - (wall << 6)) : ((wall << 6) - ori)) * inverse[abs_dir[8:0]]) >> 8;
        end
    end
end

endmodule
