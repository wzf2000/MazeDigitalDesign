module mod_top (
    // 时钟、复位
    input  wire clk_100m,           // 100M 输入时钟
    input  wire reset_n,            // 上电复位信号，低有效

    // 开关、LED 等
    input  wire clock_btn,          // 左侧微动开关，推荐作为手动时钟，带消抖电路，按下时为 1
    input  wire reset_btn,          // 右侧微动开关，推荐作为手动复位，带消抖电路，按下时为 1
    input  wire [3:0]  touch_btn,   // 四个按钮开关，按下时为 0
    input  wire [15:0] dip_sw,      // 16 位拨码开关，拨到 “ON” 时为 0
    output wire [31:0] leds,        // 32 位 LED 灯，输出 1 时点亮
    output wire [7: 0] dpy_digit,   // 七段数码管笔段信号
    output wire [7: 0] dpy_segment, // 七段数码管位扫描信号

    // PS/2 键盘、鼠标接口
    input  wire        ps2_clock,   // PS/2 时钟信号
    input  wire        ps2_data,    // PS/2 数据信号

    // // USB 转 TTL 调试串口
    // output wire        uart_txd,    // 串口发送数据
    // input  wire        uart_rxd,    // 串口接收数据

    // 4MB SRAM 内存
    inout  wire [31:0] base_ram_data,   // SRAM 数据
    output wire [19:0] base_ram_addr,   // SRAM 地址
    output wire [3: 0] base_ram_be_n,   // SRAM 字节使能，低有效。如果不使用字节使能，请保持为0
    output wire        base_ram_ce_n,   // SRAM 片选，低有效
    output wire        base_ram_oe_n,   // SRAM 读使能，低有效
    output wire        base_ram_we_n,   // SRAM 写使能，低有效

    // HDMI 图像输出
    output wire [7: 0] video_red,   // 红色像素，8位
    output wire [7: 0] video_green, // 绿色像素，8位
    output wire [7: 0] video_blue,  // 蓝色像素，8位
    output wire        video_hsync, // 行同步（水平同步）信号
    output wire        video_vsync, // 场同步（垂直同步）信号
    output wire        video_clk,   // 像素时钟输出
    output wire        video_de     // 行数据有效信号，用于区分消隐区

    // // RS-232 串口
    // input  wire        rs232_rxd,   // 接收数据
    // output wire        rs232_txd,   // 发送数据
    // input  wire        rs232_cts,   // Clear-To-Send 控制信号
    // output wire        rs232_rts,   // Request-To-Send 控制信号

    // // SD 卡（SPI 模式）
    // output wire        sd_sclk,     // SPI 时钟
    // output wire        sd_mosi,
    // input  wire        sd_miso,
    // output wire        sd_cs,       // SPI 片选，低有效
    // input  wire        sd_cd,       // 卡插入检测，0 表示有卡插入
    // input  wire        sd_wp,       // 写保护检测，0 表示写保护状态

    // // SDRAM 内存，信号具体含义请参考数据手册
    // output wire [12:0] sdram_addr,
    // output wire [1: 0] sdram_bank,
    // output wire        sdram_cas_n,
    // output wire        sdram_ce_n,
    // output wire        sdram_cke,
    // output wire        sdram_clk,
    // output wire [15:0] sdram_dq,
    // output wire        sdram_dqmh,
    // output wire        sdram_dqml,
    // output wire        sdram_ras_n,
    // output wire        sdram_we_n,

    // // GMII 以太网接口、MDIO 接口，信号具体含义请参考数据手册
    // output wire        eth_gtx_clk,
    // output wire        eth_rst_n,
    // input  wire        eth_rx_clk,
    // input  wire        eth_rx_dv,
    // input  wire        eth_rx_er,
    // input  wire [7: 0] eth_rxd,
    // output wire        eth_tx_clk,
    // output wire        eth_tx_en,
    // output wire        eth_tx_er,
    // output wire [7: 0] eth_txd,
    // input  wire        eth_col,
    // input  wire        eth_crs,
    // output wire        eth_mdc,
    // inout  wire        eth_mdio
);

/* =========== Demo code begin =========== */
wire clk_in = clk_100m;

// PLL 分频演示，从输入产生不同频率的时钟
wire clk_vga;
wire clk_ps2;
ip_pll u_ip_pll(
    .inclk0 (clk_in  ),
    .c0     (clk_vga ),  // 25MHz 像素时钟
    .c1     (clk_ps2)
);

// 七段数码管扫描演示
reg [31: 0] number;
dpy_scan u_dpy_scan (
    .clk     (clk_in      ),
    .number  (number      ),
    .dp      (7'b0        ),
    .digit   (dpy_digit   ),
    .segment (dpy_segment )
);

// 自增计数器，用于数码管演示
reg [31: 0] counter;
always @(posedge clk_in or posedge reset_btn) begin
    if (reset_btn) begin
	     counter <= 32'b0;
		  number <= 32'b0;
	 end else begin
        counter <= counter + 32'b1;
        if (counter == 32'd5_000_000) begin
            counter <= 32'b0;
            number <= number + 32'b1;
        end
	 end
end

// 图像输出演示，分辨率 800x600@75Hz，像素时钟为 50MHz，显示渐变色彩条
wire [11:0] hdata;  // 当前横坐标
wire [11:0] vdata;  // 当前纵坐标

// 生成彩条数据，分别取坐标低位作为 RGB 值
// 警告：该图像生成方式仅供演示，请勿使用横纵坐标驱动大量逻辑！！
// assign video_red = vdata < 200 ? hdata[8:1] : 0;
// assign video_green = vdata >= 200 && vdata < 400 ? hdata[8:1] : 0;
// assign video_blue = vdata >= 400 ? hdata[8:1] : 0;

localparam [0:7499][23:0] start_img = {
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011111110111111101111,
       24'b101111011011111010111110,
       24'b110100001100111111001111,
       24'b111011111110101111101011,
       24'b111011011110101011101000,
       24'b111101101111010011110010,
       24'b111110101111100111110111,
       24'b110010111100101111001011,
       24'b110000011100001011000010,
       24'b110001101100011011000110,
       24'b101111111011111110111111,
       24'b111010101110101011101010,
       24'b110111001101110011011100,
       24'b101101111011011110110111,
       24'b101100101011001110110101,
       24'b111011011110110111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100101111001011110010,
       24'b110000111100001111000011,
       24'b110000101100001011000010,
       24'b111000001110000111100001,
       24'b111101111111011111110111,
       24'b101011111011000010110011,
       24'b111001011110010111100011,
       24'b111110101111100011110011,
       24'b101110111011111010111111,
       24'b101100011011001110110100,
       24'b110000111100001111000011,
       24'b110000101100001111000011,
       24'b101111101011111110111111,
       24'b110001101100011011000110,
       24'b110010001100100011001000,
       24'b110001111100011111000111,
       24'b101111011011110110111101,
       24'b111010001110100011101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111111011111110111111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001010100010100100100101,
       24'b001001110010011000100011,
       24'b001001010010001100011111,
       24'b001010000010010100100010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100111111001111110011111,
       24'b010101000101010001010110,
       24'b000000000000000000000000,
       24'b000101000000111100001010,
       24'b111000001101110111011001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011011100110111001101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001011110010111000101110,
       24'b110100101101000111010000,
       24'b001100010010111100101101,
       24'b011001000101111101010111,
       24'b101000111001100110001011,
       24'b010111110101100101010001,
       24'b001010000010010100100100,
       24'b000000000000000000000000,
       24'b001101100011010100110001,
       24'b010000100100000000111011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100001101000011010000110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110000001100000011000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100011011000110110001110,
       24'b101011001010100110100110,
       24'b011101110111000001101000,
       24'b100111101001001010000011,
       24'b111100001110110011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100001101000011010000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b011000010101110101011001,
       24'b111110011111100011110110,
       24'b100101011000111010000101,
       24'b001101110011001000101101,
       24'b010000110100000000111100,
       24'b011011010110100001100010,
       24'b100010001000010001111001,
       24'b010000000011111100111000,
       24'b010000100100000000111010,
       24'b001010100010011100100100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b011111100111111001111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001001100010011000100,
       24'b000010010000100100001001,
       24'b000011000000110000001100,
       24'b000100110001010000010100,
       24'b000010010000100100001001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100000001000000001111,
       24'b000011110000111100010000,
       24'b000001000000010000000100,
       24'b100110101001101010011011,
       24'b111111111111111111111111,
       24'b111000001101010010111111,
       24'b110100101100010110110010,
       24'b111011011110100111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011101100111011001110,
       24'b000000000000000000000000,
       24'b001001100010010000100001,
       24'b101010011010010110011110,
       24'b110111001101101111011000,
       24'b100000010111110001110111,
       24'b000110010001011100010100,
       24'b000000000000000100000010,
       24'b000111110001111100011111,
       24'b010111000101100101010110,
       24'b010101010101001101001111,
       24'b000100000000111000001111,
       24'b000000000000000000000000,
       24'b000011110001000000001111,
       24'b000011110000111100001111,
       24'b000011110000111100001111,
       24'b000001000000010000000100,
       24'b100010001000100010001000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101111111011111110111,
       24'b111010001110100011101000,
       24'b111010101110101111101011,
       24'b111100011111001011110010,
       24'b100111101001110110011011,
       24'b000110010001011100010001,
       24'b100010111000001001111000,
       24'b101110001011000010101000,
       24'b111011011110110011101100,
       24'b111011011110110111101101,
       24'b111001001110010011100100,
       24'b111101111111011111110111,
       24'b011100110111000001101100,
       24'b001101100011010000110000,
       24'b011100100110111001100101,
       24'b111011101110110011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100111111001111110011,
       24'b000010100000101000001011,
       24'b000110100001101000010110,
       24'b011001000110001001011101,
       24'b101111101011111010111110,
       24'b001101100011001100110011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b110010011100100111001010,
       24'b111010011110100111101011,
       24'b111010011110100111101010,
       24'b111101111111011111111000,
       24'b111111001111110011111100,
       24'b111111001111110011111100,
       24'b111111101111111011111110,
       24'b111101111111011111110111,
       24'b111000111110001111100011,
       24'b111101001111010011110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010011100011011000010,
       24'b101110001010111110011101,
       24'b101101111010110010011100,
       24'b110110111101010111001111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010101110101100001011001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100110011001101110011010,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101011111010111110101,
       24'b111101101111011011110110,
       24'b111111111111111111111111,
       24'b110101011101010111010101,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b001110110011011100110110,
       24'b110010011100011111001001,
       24'b001101110011010100110011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b111000011110000111100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100101110111111101001,
       24'b101101111010111010011101,
       24'b000110010001100100010100,
       24'b010110100101100101011000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100100101001001010001,
       24'b000000110000001100000011,
       24'b000100000001000000010001,
       24'b000110010001101000011011,
       24'b001000000001111100011111,
       24'b010101000101000101001110,
       24'b010110100101011101010100,
       24'b000110010001100100011001,
       24'b000110110001101100011011,
       24'b001001000010010000100100,
       24'b000101010001010100010101,
       24'b000000000000000000000000,
       24'b000000110000001000000010,
       24'b001011100010110100101101,
       24'b110010011100100111001001,
       24'b001010010010100100101000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110100001101000011010,
       24'b001001000010010000100100,
       24'b000111000001110000011100,
       24'b000111010001110100011101,
       24'b000111000001110000011100,
       24'b000111010001110100011101,
       24'b000100010001000100010010,
       24'b011011100110110101101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010111110100111100010,
       24'b001100010010111000101000,
       24'b000000000000000000000000,
       24'b100010011000010110000001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010010100100101001001011,
       24'b000000000000000000000000,
       24'b000100010001000100010001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000100000001000000010,
       24'b000000000000000000000000,
       24'b001010100010101000101010,
       24'b110101111101011111010111,
       24'b000111100001111000011111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100100011000111110001100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100100011001000010001110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010110110101100101011001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100110101001101010011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000100000001000000010000,
       24'b000000000000000000000000,
       24'b001001010010010100100101,
       24'b110100001101000011010000,
       24'b000111100001111000011110,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001010000010011000011101,
       24'b111011001110100011011110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100101101001011010010111,
       24'b000000000000000000000000,
       24'b000000110000001100000010,
       24'b010111100101101101011011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010001100100011001000110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b011110010111100101111001,
       24'b110000111100001111000011,
       24'b101110011011100110111001,
       24'b101110011011100110111001,
       24'b101110011011100110111001,
       24'b101110101011101010111010,
       24'b110000001100000011000000,
       24'b100110111001101110011011,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000111110001111100011111,
       24'b110011101100111011001110,
       24'b001000000010000100100001,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b101000111010001110100011,
       24'b110001011100010111000101,
       24'b110000001100000011000000,
       24'b110000001100000011000000,
       24'b110000001100000011000000,
       24'b101101111011100010111001,
       24'b110101001101001011001110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101101111011111111001,
       24'b111111111111111111111111,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111110111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001011010010110100101,
       24'b000000000000000000000000,
       24'b000101110001001100001111,
       24'b110011001100100011000001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100000101000001010000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101110111011101110111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011101110111011101110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000010010000100100001,
       24'b110011111100111111001111,
       24'b001000000010000000100000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110101111101111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011111110111011101101,
       24'b010110100101100001010100,
       24'b000111010010000000100010,
       24'b010111010101110001011001,
       24'b101001001001111110010110,
       24'b010010100100100101001010,
       24'b001111100011111100111110,
       24'b010001010100010101000100,
       24'b010111100101111001011110,
       24'b010011110100111101010000,
       24'b010110110101101001010111,
       24'b011101110111010001110010,
       24'b100110001001000010001011,
       24'b011001100110001101100001,
       24'b010010010100101001001010,
       24'b010000010100000101000001,
       24'b010111110101111001011011,
       24'b100001001000000001111011,
       24'b001111110011111101000000,
       24'b011010000110100001100101,
       24'b101100011010110010100110,
       24'b110001101011111010110101,
       24'b110000011011110010110010,
       24'b110011001100100010111110,
       24'b011001010110001101011110,
       24'b010001110100100001000111,
       24'b010001010100010001000100,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010000010100000101000001,
       24'b010110110101101101011011,
       24'b001100110011001100110011,
       24'b000000000000000000000000,
       24'b000000100000000100000001,
       24'b010110000101011101010111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010011100100111001001110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100111111001111110011111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100011101000111010001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000010010000100100001,
       24'b110011111100111111001111,
       24'b001000000010000000100000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001101000011010000110100,
       24'b010010000100100001001000,
       24'b010001010100010101000110,
       24'b010001010100010101000100,
       24'b011011000110101001101001,
       24'b100100011000111010001100,
       24'b100100011000110110001001,
       24'b011010100110011001100011,
       24'b101000111010000010011001,
       24'b100010001000011010000001,
       24'b010011000100110001001011,
       24'b010000000100000001000001,
       24'b010011000100101101001011,
       24'b101111111011100110110010,
       24'b100000010111110001110111,
       24'b001110110011101100111011,
       24'b010010000100100001001000,
       24'b010111010101110101011101,
       24'b010100110101001101010011,
       24'b010010110100101101001011,
       24'b010000100100001001000010,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010001010100010101000101,
       24'b010001000100010001000100,
       24'b010000010100000001000000,
       24'b010000000011111000111101,
       24'b011001000110010101100001,
       24'b011000110110000001100000,
       24'b100100101000110110000110,
       24'b011001000110000001011111,
       24'b101001111010000010011000,
       24'b110110111101010111001000,
       24'b100011011000101110000010,
       24'b111000011110000111011111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100101101000111010001,
       24'b001101110011001000101100,
       24'b010001010011111100110110,
       24'b001101110011001100101110,
       24'b010010100100010100111110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010111000101100001010001,
       24'b001101100011001100101101,
       24'b100001000111110001110011,
       24'b000010010000011000000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001001010010001100100001,
       24'b101111011011000010100001,
       24'b011111110111011001101011,
       24'b100111011001011110001010,
       24'b101101011010100110011001,
       24'b110100011100001010110010,
       24'b110000101011011110100101,
       24'b100001111000000101110100,
       24'b001011010010110100101000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001111010011110100111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010000100100001001000010,
       24'b000000000000000000000000,
       24'b000010100000101000001010,
       24'b101100101011001010110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100011101000111010001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111110001111100011111,
       24'b110011111100111111001111,
       24'b000111110001111100011111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001110000010000000100,
       24'b000000010000000000000000,
       24'b001010000010001100011101,
       24'b001110000011001000101101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010000100011110100110111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010110100101001101001100,
       24'b011101010110110101100110,
       24'b010111110101101001010010,
       24'b010001110100000000111001,
       24'b000101000000111100001110,
       24'b011010010110001101011010,
       24'b011110100111001101100011,
       24'b011101100111001001101000,
       24'b111101001111001011101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010101110100111101000,
       24'b100111101001001110000111,
       24'b110000111011100110101101,
       24'b100000010111110001110110,
       24'b010010000100011101000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001100000010111100101100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101011101010010010010100,
       24'b110111101101000010111101,
       24'b110001011011011110101000,
       24'b101100101010011010010101,
       24'b100110001001000110000100,
       24'b011011010110010101011011,
       24'b000110100001011000010100,
       24'b000000010000000100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001011010010110100101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010001110100011101000111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100111001001110010011100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010101100101011001010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b110001101100011011000110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101100001001000010000,
       24'b001001110010010000100001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001011000010011100100010,
       24'b010011010100100101000011,
       24'b000110110001100100010111,
       24'b000000000000000000000000,
       24'b001100000010110100100111,
       24'b000000000000000000000000,
       24'b000001010000011000000101,
       24'b010011100100101101000110,
       24'b001011110010110000101000,
       24'b010011100100110101000100,
       24'b110011101100111111001101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111101101110111011011,
       24'b011111100111011101101111,
       24'b010010000100001100111110,
       24'b000010000000011100000110,
       24'b000000000000000000000000,
       24'b011111100111111101111111,
       24'b100100011001000110010001,
       24'b100101011001010010010100,
       24'b101011011010110110101110,
       24'b101001101010011110100111,
       24'b101000101010001110100011,
       24'b101010001010100010101001,
       24'b100000001000000110000010,
       24'b100010101000101010001011,
       24'b100011011000110110001101,
       24'b100010111000101110001011,
       24'b011111100111111101111111,
       24'b110001101100010010111101,
       24'b111011001110011111011111,
       24'b111000011101110011010111,
       24'b110111111101110011010110,
       24'b110000011100000010111001,
       24'b101110011011011010110011,
       24'b100100101001001010010010,
       24'b101000001010000110100001,
       24'b101100001011000010110000,
       24'b101001111010011110100111,
       24'b101010101010101110101011,
       24'b100100111001001110010011,
       24'b100011011000110110001101,
       24'b100100111001001110010011,
       24'b101011011010110110101101,
       24'b101011111010111110101111,
       24'b101011011010110110101101,
       24'b101011011010110110101101,
       24'b101011011010110110101101,
       24'b101000101010001010100010,
       24'b110010111100101111001011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100001101000011010000,
       24'b101000001010000010100000,
       24'b101000001010000010100000,
       24'b111100011111000111110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101010001010100010101000,
       24'b101001001010010010100101,
       24'b101101101011011010110110,
       24'b111111111111111111111111,
       24'b101110001011100010111000,
       24'b101001101010011010100110,
       24'b110000101011111110111101,
       24'b101110111011100110110111,
       24'b101011111010111110101111,
       24'b101011011010110110101101,
       24'b101011001010110010101100,
       24'b101010001010100110101001,
       24'b101111101011111010111110,
       24'b101111101011111010111110,
       24'b101011001010110110101101,
       24'b101110011011100110111001,
       24'b101000101010001010100010,
       24'b100011001000110010001100,
       24'b100101011001010110010101,
       24'b101011011010110110101101,
       24'b101010111010101110101011,
       24'b101011001010110010101100,
       24'b101011101010111010101110,
       24'b101001011010011010100110,
       24'b101010001010100110101001,
       24'b101010111010101010101011,
       24'b101110001011100010111001,
       24'b101100011011000110110001,
       24'b101011111010111110101111,
       24'b101001101010011110100111,
       24'b100101101001100010011001,
       24'b101010111010110010101100,
       24'b110010101100100111001001,
       24'b101101101011011110110111,
       24'b100001001000011010001001,
       24'b100000101000010010000111,
       24'b110100111101001111010011,
       24'b110001001100010011000100,
       24'b011010000110001101011100,
       24'b101101111010111010011111,
       24'b101100101010100110011101,
       24'b100111111001100010001000,
       24'b111011101110110011100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111101101110111011100,
       24'b000110100001101000011010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010010000100100001010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111101101111011011100,
       24'b111001111110011111100111,
       24'b111011001110110011101101,
       24'b110111111110000011100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101101101011111011001,
       24'b111000111110010011100110,
       24'b111111111111111111111111,
       24'b111100001110111111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100011111000111110001,
       24'b111010101110101011101010,
       24'b111011001110110111101101,
       24'b111100011111000111110001,
       24'b111100101111001011110010,
       24'b111100101111001011110010,
       24'b111001101110011011100110,
       24'b110010011100100111001001,
       24'b110010011100100111001001,
       24'b110010011100100111001001,
       24'b110010011100100111001001,
       24'b111000111110001111100011,
       24'b111100101111001011110010,
       24'b111100101111001011110010,
       24'b110101111101011111010111,
       24'b110010011100100111001001,
       24'b110000101100001011000010,
       24'b110011111100111111001111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b110010011100100111001001,
       24'b111011111111000011110000,
       24'b111100001111000011110000,
       24'b111101001111010011110011,
       24'b110100111101010011010100,
       24'b111011001110110011101100,
       24'b111100101111001011110010,
       24'b111010011110101011101010,
       24'b111010011110101011101010,
       24'b111010001110100011101000,
       24'b111010101110101011101010,
       24'b111100001111000011110000,
       24'b111100101111001011110010,
       24'b111011011110110111101101,
       24'b111010111110101111101011,
       24'b111011111110111111101111,
       24'b111000001110001011100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111001001110010011100101,
       24'b111011101110111111101111,
       24'b111010011110100111101001,
       24'b110101001101010111010110,
       24'b111110101111100011111001,
       24'b111111001111101011111010,
       24'b111101001111010011110100,
       24'b111100101111001111110010,
       24'b111011111110111111101111,
       24'b111010111110101111101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111100111111000,
       24'b110101111101101111011100,
       24'b110110111101111011011111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101111111011011110011,
       24'b101110001011100110111001,
       24'b100010011000000101110111,
       24'b101000011001101010010001,
       24'b100110111001011010001101,
       24'b011000110101111101010110,
       24'b110011001100110011001000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111111101111111011111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001110000011100000111,
       24'b111001011110010111100101,
       24'b111111111111111111111111,
       24'b101100101011010010110110,
       24'b010000100100001100111100,
       24'b001011110010110100101001,
       24'b000000000000000000000000,
       24'b000001000000010100000101,
       24'b101010001010011110100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011011100110111001101100,
       24'b000010000000011100000100,
       24'b000000000000000000000000,
       24'b000000110000001100000010,
       24'b000111110001110000011000,
       24'b111010001110100011101000,
       24'b111111111111111111111111,
       24'b110001111100100011001000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101110001011100010111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100000101000001010000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010110000101000000110,
       24'b000011100000110000000111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100010001000100010001,
       24'b000100000001000000010000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100000011000000010000000,
       24'b111111111111111111111111,
       24'b110001111100011111000111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001011010010101100101001,
       24'b010010010100010001000010,
       24'b001011110010110000101010,
       24'b000101110001100100010111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000011110000111000001100,
       24'b101110101011000110100110,
       24'b010000110100000000111100,
       24'b000100010001000100001110,
       24'b011100100110111101101000,
       24'b100101001000101101111110,
       24'b110100111100100110111001,
       24'b011110000111001001101010,
       24'b001100110011000000101101,
       24'b011000110110000001011100,
       24'b000101000001001100010011,
       24'b000100100001000100010000,
       24'b000000000000000000000000,
       24'b101110001011100110111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000100000001000000010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001110000011100000111,
       24'b111001001110010011100101,
       24'b111111111111111111111111,
       24'b101111101011111010111101,
       24'b010110100101100001001110,
       24'b001001010010001000011111,
       24'b000000000000000000000000,
       24'b011111000111011101101101,
       24'b001001010010001000100001,
       24'b100001011000011010001000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110111001100110011001,
       24'b100011101000011101111011,
       24'b111011011110001011001110,
       24'b001100110011000100101011,
       24'b000000000000000000000000,
       24'b001000010001111000011100,
       24'b111101111111100011111000,
       24'b111111111111111111111111,
       24'b101111001011110010111100,
       24'b000000000000000000000000,
       24'b000000100000000100000001,
       24'b001110010011010000110001,
       24'b000101110001010000010010,
       24'b000101100001011000010110,
       24'b000001000000010000000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110000001100000011000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010001110100011101000111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111100001110100011001,
       24'b010010010100011101000000,
       24'b000011110000111100001110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100000001000000010000,
       24'b000001000000010000000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100000101000001010000010,
       24'b111111111111111111111111,
       24'b110101111101010011010001,
       24'b001111100011101000110101,
       24'b000111010001110000011010,
       24'b010110100101011101010001,
       24'b100100011000100101111111,
       24'b001010000010011000100100,
       24'b000000000000000000000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010111110101101001010101,
       24'b000010010000011100000111,
       24'b000101010001001100001111,
       24'b000101110001011000010100,
       24'b011101110111000001101011,
       24'b100000100111010101101011,
       24'b011000000101101001010110,
       24'b011111010111011101110000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101111101011111010111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010000000100000001000,
       24'b111001011110010111100100,
       24'b111111111111111111111111,
       24'b111111011111110111111011,
       24'b011110110111011001101000,
       24'b000000000000000000000000,
       24'b010010110100010101000011,
       24'b101110001010111110100011,
       24'b011001000101111101010111,
       24'b010100100100110101001000,
       24'b111000001101111011011100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101101111010011110001,
       24'b001111100011100000101110,
       24'b010110110101010001001110,
       24'b100110011001000110000101,
       24'b110100111100101110111100,
       24'b001010110010101000100111,
       24'b000000000000000000000000,
       24'b111000101110000111100010,
       24'b111111111111111111111111,
       24'b110100011100111111010000,
       24'b000111000001101000011010,
       24'b000000100000001000000010,
       24'b001011100010110100101100,
       24'b000110000001011100010110,
       24'b000101010001010100010101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b001000100010001000100010,
       24'b111111101111111011111110,
       24'b111111111111111111111111,
       24'b110011011100100010111111,
       24'b001110100011010000101100,
       24'b000000000000000000000000,
       24'b000111010001101100011000,
       24'b100001000111111101110110,
       24'b000001000000010000000011,
       24'b001000110001111100011101,
       24'b010001010100001000111110,
       24'b000100110001000000001110,
       24'b000000000000000000000000,
       24'b000011000000110000001100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100000001000000110000001,
       24'b111111111111111111111111,
       24'b101101001011010110110100,
       24'b000000000000000000000000,
       24'b000111110001111100011110,
       24'b011010000110001001011100,
       24'b101010011010001010010110,
       24'b011001000101110101010101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010100110100111001000111,
       24'b101010011010001010011001,
       24'b001000100001111000011100,
       24'b011111010111011001101110,
       24'b011001000101111101010111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101110001011100010111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101110111011101,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001000000010000000100,
       24'b111000101110001011100010,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b101000001001011110001100,
       24'b000010100000101000001010,
       24'b010111100101101001010100,
       24'b001110100011010100110110,
       24'b011001000110001001011011,
       24'b001110110011011000110010,
       24'b001001010010001000100000,
       24'b111000011110000111100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010001100100111001100,
       24'b100011101000100101111110,
       24'b011001010110000101010111,
       24'b000000000000000000000000,
       24'b001101010011001100110001,
       24'b111000101101010111001000,
       24'b001110110011100100110111,
       24'b000000000000000000000000,
       24'b110110101101100111011001,
       24'b111111111111111111111111,
       24'b110011101100110111001101,
       24'b000110000001011000010110,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001100000011000000110,
       24'b000100000001000000010000,
       24'b000100010001000100010001,
       24'b000100100001001000010010,
       24'b000100010001000100010001,
       24'b000100100001001000010010,
       24'b000100010001000100010001,
       24'b000100010001000100010001,
       24'b000101100001011000010110,
       24'b000011010000111000001110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000100010001000100010,
       24'b111111101111111011111110,
       24'b111111111111111111111111,
       24'b110101001100111111001000,
       24'b010100000100101101000110,
       24'b000011010000110100001101,
       24'b010110110101011101010001,
       24'b101001001001110010001111,
       24'b001001110010011100100110,
       24'b101100111010110010011111,
       24'b101001001010000110010100,
       24'b010100110101000001001110,
       24'b000110010001100000011001,
       24'b001111110011111100111111,
       24'b001111000011110000111100,
       24'b000000100000001000000010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100000101000001010000010,
       24'b111111111111111111111111,
       24'b110010101100101111001011,
       24'b000110100001100000010110,
       24'b000000000000000000000000,
       24'b000010000000011100000111,
       24'b010001010100010000111110,
       24'b101000111001110010001111,
       24'b000100100001001000010010,
       24'b000011100000111000001110,
       24'b000011100000111000001110,
       24'b010001000100001000111101,
       24'b101010111010010110011010,
       24'b010111110101101001010101,
       24'b001011000010101100101011,
       24'b001010000010011100100111,
       24'b001100110011000000110001,
       24'b100010101000011001111110,
       24'b011110010111010001101101,
       24'b001100010011000000110001,
       24'b100010101000011001111101,
       24'b011101000111000101101010,
       24'b000011100000111100001111,
       24'b000100010001000100010001,
       24'b000011110000111100001111,
       24'b000011000000110000001100,
       24'b110000101100001011000010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100100001001000010010,
       24'b111010011110100111101001,
       24'b111111111111111111111111,
       24'b110100011100111111001101,
       24'b000010010000011100000110,
       24'b000000000000000000000000,
       24'b000100000001000000001110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000010010000100100001,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011001110110011101010,
       24'b101000101001110010010011,
       24'b010111000101010101001101,
       24'b000010010000100000001001,
       24'b000000000000000000000000,
       24'b001001110010010000100101,
       24'b001011100010011100100100,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b110111001101110011011100,
       24'b111111111111111111111111,
       24'b110000011100000111000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110100001101000011010,
       24'b111011001110110011101100,
       24'b111100111111001111110011,
       24'b111011111110111111101111,
       24'b111100001111000011110000,
       24'b111011111110111111101111,
       24'b111100001111000011110000,
       24'b111100001111000011110000,
       24'b111011111110111111101111,
       24'b111101101111011011110110,
       24'b101001001010001110100011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000110010001100100011,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111001011110010111100100,
       24'b111000001110000111100010,
       24'b111011011110110111101100,
       24'b111101101111011011110111,
       24'b111110001111100011111000,
       24'b111110011111101011111000,
       24'b111110001111100011110110,
       24'b111001111110011011100110,
       24'b111101001111010011110011,
       24'b111111001111110011111100,
       24'b111101111111011111110111,
       24'b010101100101011001010110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010010100100101101001010,
       24'b111010101110100111101001,
       24'b111111111111111111111111,
       24'b111001001110001011100000,
       24'b101101111010111010011110,
       24'b001010100010011100100001,
       24'b000000000000000000000000,
       24'b001010100010011000100100,
       24'b111000111110000111100001,
       24'b111100111111001011110011,
       24'b111011011110110111101101,
       24'b111011011110110011101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011111110111111101101,
       24'b111111111111111111111111,
       24'b111110101111100111111001,
       24'b111010111110101111101100,
       24'b111001101110011011100101,
       24'b111101001111010011110010,
       24'b111101011111011011110101,
       24'b111010001110100011100110,
       24'b111101111111011111110110,
       24'b111011011110111011101110,
       24'b111100001111000011110000,
       24'b111011111110111111101111,
       24'b111010101110101011101010,
       24'b111110111111101111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101010001010100010110,
       24'b111101011111010111110101,
       24'b111111111111111111111111,
       24'b110001111100011111001010,
       24'b000000000000000000000000,
       24'b000010110000100000000111,
       24'b000100010000111100001111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001100000011100000111,
       24'b000011000000110100001101,
       24'b000000000000000000000000,
       24'b010000100100001001000011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110110111100101110001,
       24'b011100000110100001011100,
       24'b010111010101011101010000,
       24'b010111000101011001001111,
       24'b000100110001001000010001,
       24'b000101010001001100010010,
       24'b010001010100010001000011,
       24'b000000000000000000000000,
       24'b000000100000001000000010,
       24'b110110111101101111011011,
       24'b111111111111111111111111,
       24'b110000111100001111000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111010001110100011101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110000101100000111000000,
       24'b000000000000000000000000,
       24'b000110000001011000010111,
       24'b000000000000000000000000,
       24'b000111100001111100011111,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010101000101010001010100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b011010100110101001101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001111100100011000111,
       24'b101000111001101010001011,
       24'b010110010101010101001100,
       24'b000000100000000100000010,
       24'b011011100110100101100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110001101100011011000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001010000010100100101000,
       24'b010100000101000001001110,
       24'b111000101110000111100000,
       24'b111111111111111111111111,
       24'b111001101110011111100011,
       24'b100100001000100001111001,
       24'b110010111011111110110000,
       24'b010110100101010101010000,
       24'b000101100001011100010111,
       24'b001011000010110000101100,
       24'b000000000000000000000000,
       24'b000001010000010100000101,
       24'b000001000000001100000011,
       24'b000000000000000000000000,
       24'b100101101001011010010110,
       24'b110010111100100011000001,
       24'b010011000100011100111101,
       24'b000110110001101100011001,
       24'b001010100010101000101010,
       24'b010101110101000101001100,
       24'b010001100100010101000010,
       24'b010010110100101101001000,
       24'b010010100100100001000110,
       24'b000000000000000000000000,
       24'b000000100000001000000010,
       24'b110111001101110011011100,
       24'b111111111111111111111111,
       24'b110001001100010011000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111100001111000011110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010011100100011001000,
       24'b000001110000010000000011,
       24'b000010100000100100001001,
       24'b000000000000000000000000,
       24'b000111100001111100011111,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101110111011101,
       24'b001001010010010100100101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100100011001000110010001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110111101101111011010,
       24'b110000011011100110101010,
       24'b011100010110111001100101,
       24'b000000000000000000000000,
       24'b010011100100101101000111,
       24'b111011001110101111101000,
       24'b110110001101011111010110,
       24'b110001101100011011000111,
       24'b110011101100111111001111,
       24'b110101111101100011011000,
       24'b101110101011101010111100,
       24'b110101001101010011010100,
       24'b110011111100111011001100,
       24'b111001111110011011100100,
       24'b111100101111000011101110,
       24'b111100001111000011110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000001110000011100000,
       24'b000011100000101100001101,
       24'b000000000000000000000000,
       24'b000110100001101000011001,
       24'b010010010100011101000011,
       24'b111001011110010011100011,
       24'b111111111111111111111111,
       24'b111111011111101011110110,
       24'b111011111110010111010010,
       24'b111011101110010111010011,
       24'b000110110001100000010101,
       24'b001000110010001100100101,
       24'b111000111110010011100100,
       24'b001001100010011000100110,
       24'b000000100000001000000010,
       24'b000111010001101100011010,
       24'b001111000011100100110110,
       24'b000011100000101100001001,
       24'b010110110101010101001111,
       24'b001100110010111100101011,
       24'b000001010000011100001000,
       24'b000000000000000000000000,
       24'b010010000100011101001000,
       24'b111010011110100011101000,
       24'b000101000001010000010100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b110111001101110011011100,
       24'b111111111111111111111111,
       24'b110001011100010011000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111000001110000011100,
       24'b111101101111011011110110,
       24'b111111001111110011111100,
       24'b111110101111101011111010,
       24'b111101101111011111110111,
       24'b111111001111101111111011,
       24'b111111111111111111111111,
       24'b111100011111001011110010,
       24'b111100101111000011110001,
       24'b111110101111101011111010,
       24'b101000101010001110100010,
       24'b010011010100100101000001,
       24'b010010010100011101000011,
       24'b000000000000000100000010,
       24'b000000100000001000000011,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110001011100010111000,
       24'b000011010000110100001101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101011011010110110101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110111011100110111010,
       24'b100101111000111110000100,
       24'b010011000100100001000010,
       24'b000000000000000000000000,
       24'b010000010011111000111000,
       24'b111000011101011111000111,
       24'b101111101011010010100101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101110001010000010001,
       24'b011001110110000001011000,
       24'b001111000011100100110101,
       24'b001011010010101100101000,
       24'b001010000010001100011110,
       24'b001100110010110100100111,
       24'b110001111100100011001000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010100110011101100001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b111000101110010011100101,
       24'b111111111111111111111111,
       24'b110101011101001111010100,
       24'b101010101010001010010101,
       24'b100100101000101101111100,
       24'b000000000000000000000000,
       24'b000100100001001100010110,
       24'b111111111111111111111111,
       24'b111011111110111011101110,
       24'b000100100001000000001111,
       24'b000001010000010000000011,
       24'b000101010001010000010100,
       24'b000000000000000000000000,
       24'b000000010000001000000010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001010000011000000110,
       24'b111010111110110011101100,
       24'b111111111111111111111111,
       24'b000000010000000000000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b110111001101110011011100,
       24'b111111111111111111111111,
       24'b110001011100010111000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001000000010000000100,
       24'b000111100001111000011110,
       24'b001000010010000100100001,
       24'b000101110001011100010111,
       24'b000101100001011000010110,
       24'b001000100010001000100001,
       24'b101010011010010010011101,
       24'b111001001101100011001010,
       24'b011110000111001101101000,
       24'b001000010010000100100001,
       24'b000010110000101100001011,
       24'b011101000111000101101001,
       24'b010100110101000101001100,
       24'b000000000000000000000000,
       24'b010110010101010101010010,
       24'b111111101111110111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101000001010000010100000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000100000001000000010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110110001101100011011,
       24'b110001111100011111000111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011001100101111001011,
       24'b100010111000001101110111,
       24'b000111100001101100011010,
       24'b000000000000000000000000,
       24'b000101100001010000010010,
       24'b011100100110110101100110,
       24'b101101001010111010011110,
       24'b010110000101011001001111,
       24'b000000000000000000000000,
       24'b000000010000000000000000,
       24'b100000000111100001101111,
       24'b001011010010110000101011,
       24'b000111110001111100011111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b110110011101100111011000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111101011111001,
       24'b011010100110100001011111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010010000100000001000,
       24'b111001001110010111100101,
       24'b111111111111111111111111,
       24'b110010011100101111001100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000100000001100000011,
       24'b001000100010001100100011,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b100101111001011110010110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b110000001100000111000001,
       24'b111111111111111111111111,
       24'b110111101101111111011111,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b110111001101110011011100,
       24'b111111111111111111111111,
       24'b110000111100010011000100,
       24'b000000000000000000000000,
       24'b001100110011000100101111,
       24'b010010010100011101000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010010000100001000111011,
       24'b101001101001110010001111,
       24'b010000010011111000110110,
       24'b000000000000000000000000,
       24'b000010000000011100000110,
       24'b110101111101000011000011,
       24'b001010110010100000100101,
       24'b001101110011001000101100,
       24'b111010111110001011010100,
       24'b111110011111100111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100110111001101110011,
       24'b000000000000000000000000,
       24'b000100010001000100010001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001101110011011100110111,
       24'b111011001110110011101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001011100010011000011,
       24'b010100010100110101000111,
       24'b001010000010011000100101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100100001000100001101,
       24'b010011000100100101000010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b110101101101011011010110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111001011110010111100100,
       24'b001011010010100100100110,
       24'b000101000001001000010000,
       24'b000000000000000000000000,
       24'b000001010000011000000110,
       24'b111001001110010011100100,
       24'b111111111111111111111111,
       24'b111110101111101111110111,
       24'b010001110100010000111101,
       24'b000111100001110100011101,
       24'b000100010000111100001101,
       24'b001000000001111100011110,
       24'b111110011111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110110111101101111011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100011101000111010001110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000001110000011100000,
       24'b000001000000010000000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000100000001000000010,
       24'b110110111101101111011011,
       24'b111111111111111111111111,
       24'b101111011011110110111110,
       24'b000000010000000100000000,
       24'b011000100101111101011001,
       24'b001101000011000100101111,
       24'b000001000000010000000101,
       24'b000011110001000000001101,
       24'b000000000000000000000000,
       24'b001000110010001100100011,
       24'b000010000000100000001000,
       24'b000000000000000000000000,
       24'b000000100000000100000000,
       24'b001011000010101000100111,
       24'b010111100101101001010100,
       24'b000000000000000000000000,
       24'b001010100010100000100101,
       24'b110010111100001010110011,
       24'b100010111000010101111101,
       24'b011000010101110101010010,
       24'b010001000011111100111110,
       24'b111101001111010111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110100101101001011010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010110010101100101011001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110011011100010110110,
       24'b000000000000000000000000,
       24'b000110110001100100011000,
       24'b000000000000000000000000,
       24'b000000100000001000000010,
       24'b000100010001000100010001,
       24'b000101110001011100010111,
       24'b000100010001001000010000,
       24'b000100000001001000010011,
       24'b000100000001000100010010,
       24'b000011000000110000001101,
       24'b000100000001000000010000,
       24'b000100100001001000010010,
       24'b000011110000111100001111,
       24'b000100110001001000010010,
       24'b110110101101101011011011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101001101011011010111,
       24'b000100000000111000001111,
       24'b100000000111100101110010,
       24'b000100110001000100010000,
       24'b000000000000000000000000,
       24'b111001001110010011100101,
       24'b111111111111111111111111,
       24'b110011111100111111001110,
       24'b001001000010001100100000,
       24'b010001010100001100111111,
       24'b000101010001001100010001,
       24'b000011110000111000001110,
       24'b111110011111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100010101000101010001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b011010110110101101101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001010000010100000101,
       24'b110111101101111011011110,
       24'b111111111111111111111111,
       24'b101111111011111010111110,
       24'b000001100000010100000011,
       24'b010100010100110101001000,
       24'b000111110001101100011000,
       24'b000101110001010100010011,
       24'b001110000011100100110101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001010110010100100100110,
       24'b011000010101110101011000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101011101010010010011001,
       24'b101101001010101110011101,
       24'b011010010110000101011001,
       24'b011011010110101001100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010101110101011101010,
       24'b001010100010101000101011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001000000010000000011,
       24'b000011010000110000001011,
       24'b000000000000000000000000,
       24'b011110010111100101111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111111011111010111110,
       24'b000011000000101100001010,
       24'b000001010000010000000100,
       24'b000000000000000000000000,
       24'b000100110001001100010011,
       24'b111000101110000111100010,
       24'b111100001111000111110000,
       24'b111010011110101011101010,
       24'b111011011110111111110000,
       24'b111011111110111111110000,
       24'b111100001110111111101111,
       24'b111011111110111111101111,
       24'b111011111110111111101111,
       24'b111011011110110111101101,
       24'b111011011110110111101101,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111111111111,
       24'b111111101111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111101101111011011110,
       24'b000001000000010000000100,
       24'b010011110100110001001000,
       24'b001010000010010100100100,
       24'b000111100001111100011111,
       24'b111000011110000111100001,
       24'b111111111111111111111111,
       24'b110010001100100011001000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111010001110100011101,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b000011110000111100001111,
       24'b001000110010001100100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001000000010000000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100010001000100010001,
       24'b111010101110101011101010,
       24'b111111111111111111111111,
       24'b110010111100101111001011,
       24'b001011010010101100101000,
       24'b001110010011011000110011,
       24'b000111010001101100011001,
       24'b001011010010101000100111,
       24'b101101111011011010110111,
       24'b101110001011100010111000,
       24'b101100111011001110110011,
       24'b101101001011001110110011,
       24'b101100111011010010110101,
       24'b101011111010111110110000,
       24'b110010101100100011000110,
       24'b110010011100100111001010,
       24'b110000001100000111000001,
       24'b011100000111000001110001,
       24'b011101110111000001101000,
       24'b101000101001110010010011,
       24'b000101010001010000010011,
       24'b001101110011010000110001,
       24'b111111101111111011111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010101100101111001011,
       24'b000110010001100000011000,
       24'b000000000000000000000000,
       24'b000101100001010100010101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111010001101100011010,
       24'b101110001011100110111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110000001100000011000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101010001010100010101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110111101110011011100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000100000001000000011,
       24'b000101010001010100010101,
       24'b111001001110010011100100,
       24'b111111111111111111111111,
       24'b110010101100101111001011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000000010000000100000,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110111101101111011011,
       24'b111001101110011011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001100000011000000110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b110111101101111011011110,
       24'b111111111111111111111111,
       24'b110001001100010111000110,
       24'b000001000000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000010010000100100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001001100011111000110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101110001011100011001,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b101110011011100110111001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010101110101001101001110,
       24'b000111010001101100011001,
       24'b000000000000000000000000,
       24'b001101110011011000110101,
       24'b101110001011010110110100,
       24'b111110001111011111110110,
       24'b111000011110000011011110,
       24'b110100011101000111010001,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110010101100101011001010,
       24'b111001111110011111100111,
       24'b111111111111111111111111,
       24'b110000001100000011000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100010001000100010001,
       24'b110001011100010111000101,
       24'b110101011101010111010101,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110100001101000011010000,
       24'b110010111100101111001011,
       24'b110010001100100011001000,
       24'b110010011100100011001000,
       24'b110100011101000111010001,
       24'b110100101101000111010010,
       24'b110111001101101111011100,
       24'b111110111111101011110111,
       24'b111111101111110011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100101111000011101101,
       24'b111011011110101111101001,
       24'b111110101111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001000000010000000100,
       24'b111001011110010111100101,
       24'b111111111111111111111111,
       24'b110001001100011011000110,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000111100001111000011110,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001100000011000000101,
       24'b110111001101110011011100,
       24'b111111111111111111111111,
       24'b110011101100110111001100,
       24'b000011010000101100001011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110010001100000010111,
       24'b111110101111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011111011000010110000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111100001111000011111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010001100100011001000110,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b000001110000011000000110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001001000010000000011111,
       24'b001100110011001000110011,
       24'b000000110000001000000010,
       24'b000010100000100000000110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100000001000000010000000,
       24'b111111111111111111111111,
       24'b110000011100000111000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001001000010001100100001,
       24'b001000010010000000011011,
       24'b001001100010010100100010,
       24'b000111100001110000011011,
       24'b000110110001100000011000,
       24'b000000010000000000000001,
       24'b010000000011111000111011,
       24'b011100000110101101100010,
       24'b010101010101000001001010,
       24'b001100110011000000101101,
       24'b100001000111110001110010,
       24'b101100101010011110011001,
       24'b101101111010110010011101,
       24'b111010101110011011100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101110111011101,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b111001001110010011100100,
       24'b111111111111111111111111,
       24'b110110101101100011011000,
       24'b000101010001001100010011,
       24'b000101100001011000010110,
       24'b000000000000000000000000,
       24'b000110110001101100011011,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000000000000000000000000,
       24'b000101100001010100010100,
       24'b010011010100101101000110,
       24'b010111010101101101010111,
       24'b110111101101111011011110,
       24'b111111111111111111111111,
       24'b111010101110100111101000,
       24'b001011100010101100101010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010101010101000101001101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011111010111110101111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001011110010111100101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010101110101011101010111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000001100000100,
       24'b000000000000000000000000,
       24'b000100110001000000001111,
       24'b000000000000000000000000,
       24'b000111000001100100011001,
       24'b001110010011011000110010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b100000001000000010000000,
       24'b111111111111111111111111,
       24'b110000011100000111000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010010000011100000111,
       24'b000011010000110000001011,
       24'b001101100011010000110011,
       24'b000111110001110000011011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000011110000110000001010,
       24'b000011110000110100001101,
       24'b001111010011110000111000,
       24'b100000100111110001110010,
       24'b101010101010001010010110,
       24'b110000111011100010101001,
       24'b110010101011110010101100,
       24'b111011111110101111100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110111101101111011011,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101100001011000010110,
       24'b111000101110001011100010,
       24'b111111111111111111111111,
       24'b110110101101100111011001,
       24'b000100000000111100001111,
       24'b000000100000001000000010,
       24'b000000000000000000000000,
       24'b000111110001111100011111,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000101110001011100010,
       24'b000001000000010000000100,
       24'b000011110000111100001110,
       24'b000110000001011100010101,
       24'b000111000001101100011001,
       24'b111001101110011011100110,
       24'b111111111111111111111111,
       24'b110010001100011111000111,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010011010100110001001010,
       24'b111111101111111011111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011111010111110101111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001110000011100000111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010011100100111001001110,
       24'b000000000000000000000000,
       24'b000100000001000000010000,
       24'b001010010010011100100100,
       24'b000001000000001100000000,
       24'b001110010011011000110010,
       24'b000111010001110000011011,
       24'b000000000000000000000000,
       24'b011001000101111001011000,
       24'b010110100101011001001111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b011111010111110101111101,
       24'b111111111111111111111111,
       24'b101111101011111010111110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000011100000110000001011,
       24'b001110110011011000110001,
       24'b011100100110101101100000,
       24'b101001101001111010010000,
       24'b101110101011000110100100,
       24'b101110111011001010100100,
       24'b100111111001010110001010,
       24'b101100101010010110011000,
       24'b101000101001011010000111,
       24'b111001111110010111100000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101110111011101,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101010001010100010101,
       24'b111000101110001011100010,
       24'b111111111111111111111111,
       24'b110001011100010111000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111100001111000011110,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101100001011100010111,
       24'b110110001101100011011000,
       24'b111111111111111111111111,
       24'b110010001100100011001001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100100001001100010011,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011111010111110101111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111000001110000011100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010111110101111101011111,
       24'b000000000000000000000001,
       24'b001110010011100100111001,
       24'b001111010011110000111001,
       24'b000010000000100000000111,
       24'b010101000101000001001100,
       24'b000100000000111100001110,
       24'b000100100001000100010001,
       24'b001000010001111100011101,
       24'b000000000000000000000000,
       24'b000010010000100000001000,
       24'b000010000000100000001000,
       24'b000010010000100100001001,
       24'b000010000000100000001000,
       24'b000010010000100100001001,
       24'b000010000000100000001000,
       24'b000010000000100000001000,
       24'b000000000000000000000000,
       24'b100010001000100010001000,
       24'b111111111111111111111111,
       24'b110000101100001011000010,
       24'b000000110000001100000011,
       24'b000001100000011000000110,
       24'b000010000000100000001000,
       24'b000010010000100100001001,
       24'b000010000000100000001000,
       24'b000010010000100100001001,
       24'b000010000000100000001000,
       24'b000010010000100100001001,
       24'b000010010000100100001001,
       24'b000010000000100000001000,
       24'b000010000000100100001001,
       24'b000010000000100000001000,
       24'b000001010000011000000111,
       24'b000001100000011000000110,
       24'b010000010011110000111001,
       24'b001101010011001000110000,
       24'b000100100000111100010001,
       24'b011100100110110001100110,
       24'b100011001000010101111011,
       24'b000011100000111100001111,
       24'b001111110011110100111011,
       24'b100101101000111110000111,
       24'b001001100010010100100001,
       24'b110011111101000011001110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001100000011000000110,
       24'b111111101111111011111110,
       24'b111111111111111111111111,
       24'b111000001110000011100000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111110001111100011111,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000101110001011100010,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000010000000100000001000,
       24'b000111110001111100011111,
       24'b111011111110111111101111,
       24'b111111111111111111111111,
       24'b110100111101001111010011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111000001110000011100,
       24'b111110111111101111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011001010110010101100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001010000010100000100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110101111101011111001,
       24'b111101001111010011110100,
       24'b111100101111001011110011,
       24'b111111001111110011111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111101111111011,
       24'b111101101111011111110111,
       24'b111111101111111011111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101111111011111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110101111101011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111101111111111111111,
       24'b111100101111001111110100,
       24'b110111101101111111100001,
       24'b111001011110011111101010,
       24'b110000001011100010101101,
       24'b100111011001010010000101,
       24'b100100101000100101111100,
       24'b101101101010110110100000,
       24'b111011011110110111100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010010000100100001001,
       24'b110000001100000011000000,
       24'b110111111101111111011111,
       24'b101010101010101010101010,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111100001111000011110,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001000000010000000100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b101111001011110010111100,
       24'b110111101101111011011110,
       24'b101100001011000110101111,
       24'b000010000000100000001000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110110001101100011011,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100011011000110110000,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101110001011100010111,
       24'b101111001011110110111111,
       24'b110100011101000011010000,
       24'b111001001110010011100100,
       24'b110101011101011111011010,
       24'b110110111101110011011110,
       24'b111010101110101011101010,
       24'b111011001110110011101100,
       24'b111000111110010011100100,
       24'b111010011110100111101001,
       24'b111011011110110111101101,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011111110111111101111,
       24'b110111011101110111011101,
       24'b110011101100111011001111,
       24'b110101011101010011010101,
       24'b111010111110101011101011,
       24'b111011011110110111101101,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111011001110110011101100,
       24'b111010001110100011101000,
       24'b111010111110101111101011,
       24'b111001011110011011100110,
       24'b111111111111111111111111,
       24'b111000101110001011100000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111101011010010101001,
       24'b100111111001010110000111,
       24'b110000011011010110101000,
       24'b101111101011000010100011,
       24'b110110011101101111010100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111010001110100011101,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000011110000111100001,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001010100010101000101001,
       24'b000111100001111100011111,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110110001101100011011,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110001101100111010101,
       24'b000111000001111000011001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001000000010000100100000,
       24'b001111000011110000111010,
       24'b010100100100111101001010,
       24'b010000110011111100111010,
       24'b010000000011111000111010,
       24'b001100010010111100101100,
       24'b000010010000100000001000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000110000010000000100,
       24'b000010110000100100001001,
       24'b001010010010010000100011,
       24'b000101110001010000010011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001101000011000100101110,
       24'b010101110101010101010000,
       24'b010010010100011101000001,
       24'b101000011001101110010000,
       24'b001001110010010100100010,
       24'b011010010110100001100011,
       24'b111011011110000011001110,
       24'b101100011010001010010100,
       24'b110110011101101111010110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001001110010011100100111,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000101110001011100010,
       24'b000001010000010100000101,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000110110001101100011011,
       24'b111110111111101111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001101100011011000101,
       24'b000001110000100000000110,
       24'b000000000000000000000000,
       24'b000001100000010100000101,
       24'b011000100101111101011000,
       24'b011110000111011001110001,
       24'b001111010011101000110110,
       24'b010001100100001000111101,
       24'b010000110100000000111100,
       24'b001001000010001000011110,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000011010000110100001101,
       24'b000010010000100100001001,
       24'b000000000000000000000000,
       24'b000000110000001100000011,
       24'b000011010000110100001101,
       24'b000010100000100100001000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000100010001000000010000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b010111010101100101010100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001001100010011000100100,
       24'b110101001100100110111001,
       24'b110101101100011110110100,
       24'b111100101111000011101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101110011011100,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000101100001011000010110,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000001110000011100000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010010000100100001010,
       24'b111111101111111011111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101000111010001110100011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001100000011100001000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000111110001101100011000,
       24'b001101100011010000110001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000010100000101000001011,
       24'b011010100110010001011110,
       24'b010101010101000001001011,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b001001010010001100011101,
       24'b100111101001011110001100,
       24'b111110011111011011110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110001101100011011000,
       24'b000000100000001000000010,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000111010001110100011101,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111111101111111011111,
       24'b000000110000001100000011,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000011000000101100001011,
       24'b001101000011000100101111,
       24'b010000000011111000111100,
       24'b111011111110111111101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100011011000110110001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000011100000111000001110,
       24'b000101110001011000011000,
       24'b000000000000000000000000,
       24'b001001110010010100100011,
       24'b010000100100000000111100,
       24'b000000000000000000000000,
       24'b000000000000000000000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000110010001011100010110,
       24'b001000100010001000100000,
       24'b000000110000001100000011,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000100000001000000010,
       24'b000000010000000100000001,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000010100000101000001010,
       24'b000011100000111000001110,
       24'b000010110000101100001011,
       24'b000100100001001000010010,
       24'b000000000000000000000000,
       24'b000100100001001000010010,
       24'b000010110000101100001011,
       24'b000000000000000000000000,
       24'b000110010001100000010111,
       24'b010001000100001000111111,
       24'b000110010001100000010110,
       24'b000000000000000000000000,
       24'b000100010001000000010001,
       24'b100000000111100101110000,
       24'b010001000011111000111000,
       24'b000000000000000000000000,
       24'b000000000000000100000001,
       24'b000000010000000100000001,
       24'b000000000000000000000000,
       24'b000000000000000000000000,
       24'b000001010000010000000011,
       24'b110010111100101011001001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101101111011011110110,
       24'b110110111101101111011011,
       24'b110110111101101111011011,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110110001101100011011000,
       24'b111000001110000011100000,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110011111100111111001,
       24'b110110111101101111011011,
       24'b110110101101101011011010,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110110001101100011011000,
       24'b111010001110011111100111,
       24'b111111111111111111111111,
       24'b111101111111010111110011,
       24'b111101101111011011110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101111111011111110111,
       24'b110110101101101011011010,
       24'b110111001101110011011100,
       24'b111001101110010111100101,
       24'b111010111110101111101011,
       24'b110101001101010111010101,
       24'b111100101111000011101101,
       24'b111111111111111111111111,
       24'b110110101101101011011011,
       24'b110111001101110011011100,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110101101101011011010111,
       24'b110100111101001111010011,
       24'b110111011101110111011101,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110110111101101111011011,
       24'b111001001110010011100100,
       24'b111001101110011011100110,
       24'b111001011110010111100101,
       24'b111010111110101111101011,
       24'b110101101101011011010110,
       24'b111001011110010111100101,
       24'b111000111110001111100011,
       24'b110101101101011111010111,
       24'b111100101111000111101111,
       24'b111111111111111111111111,
       24'b111100111111001011110000,
       24'b110101011101011011010110,
       24'b110100001101000011010000,
       24'b111000001110000011011111,
       24'b111000011110000011011110,
       24'b110110011101100111011000,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110111101101111011011110,
       24'b110110111101101011011011,
       24'b110010001100100011001001,
       24'b111011001110110011101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
};
localparam [0:7499][23:0] end_img = {
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101111111010011110110,
       24'b111010011110100011110100,
       24'b101001011001100111101100,
       24'b011111100110101111011111,
       24'b111111001111110111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111011011110101011110110,
       24'b100110001000110111100110,
       24'b111111111111111111111110,
       24'b110111011101011111110011,
       24'b001100100001111011011000,
       24'b001011110001001011010110,
       24'b000110100000000011011001,
       24'b000011100000000011010011,
       24'b110000111011100111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111011111110111011110101,
       24'b110101111101000111110011,
       24'b101011111010011011110001,
       24'b100110011000100111100111,
       24'b101000101001001011100001,
       24'b110011001100011011101001,
       24'b001101110010001111011010,
       24'b000000000000000011010010,
       24'b010110010100000111011010,
       24'b001100010001011011010100,
       24'b000011000000000011011000,
       24'b001001110000011011011011,
       24'b010001100010101011010111,
       24'b000110000000010111011001,
       24'b100110011000100111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110001111011111111001,
       24'b110011111100101111101111,
       24'b101011001010000111101101,
       24'b100010110111101011100111,
       24'b010010010011001111100000,
       24'b001100100001010011011101,
       24'b010010100011001111010100,
       24'b001001000000100011010011,
       24'b001000110000001011011010,
       24'b000011010000000011010110,
       24'b000110100000000011010011,
       24'b001000110000001111010111,
       24'b010100110011011111011010,
       24'b010101000011110011010101,
       24'b010111000100100111100000,
       24'b101110101010110111101100,
       24'b111001001101111111110010,
       24'b100001100111010011011110,
       24'b000110000000011111010111,
       24'b100010000111010111100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b110110011101011111110100,
       24'b101010001010000111101110,
       24'b100001100111011111100101,
       24'b011001110101100011100010,
       24'b010010100011000011011010,
       24'b001010100000110111010111,
       24'b000000000000000011011010,
       24'b000000000000000011011011,
       24'b000010010000000011011000,
       24'b000000100000000011010111,
       24'b000011110000000011010101,
       24'b001111100010001011010111,
       24'b010011100011010011011010,
       24'b010011000011011111100001,
       24'b011111100110110011100100,
       24'b110011011100010011101111,
       24'b111111001111110011110110,
       24'b111111001111110011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010110101010011100100,
       24'b000000000000000011010011,
       24'b001000000000000011011100,
       24'b111100011111001011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111001111110100011111001,
       24'b101111001011010111110000,
       24'b100011001000000111101000,
       24'b011010010101011111100101,
       24'b010000110010100111011111,
       24'b000111000000000011011011,
       24'b000001110000000011011001,
       24'b000000100000000011011000,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000000000000000011011011,
       24'b000011010000000011011010,
       24'b000111100000000011011001,
       24'b010001010010110011011100,
       24'b011110010110011011100010,
       24'b101000001001001111101011,
       24'b110001001011101011110000,
       24'b111011011110100011110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101010011001110011101100,
       24'b011100110110001011011100,
       24'b010111100100101111010111,
       24'b110101111101001111110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111010111110101111110111,
       24'b110010101100011011110010,
       24'b100110111001001111101010,
       24'b011101000110010111100101,
       24'b010101000100000111100000,
       24'b001010100000110011011101,
       24'b000011010000000011011000,
       24'b000000000000000011010111,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011010111,
       24'b001010000000100011011011,
       24'b010100010011100011011111,
       24'b010100100011111111100010,
       24'b100001100111100111100111,
       24'b101111111011100011101111,
       24'b111000111110000111110101,
       24'b111101101111010111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011001110110011110001,
       24'b011011000101010111011011,
       24'b001100110010111011010110,
       24'b101010011001111011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b111100101111001111111000,
       24'b101110011011010111110001,
       24'b101000011001011111101011,
       24'b100101101000100011100101,
       24'b010101000100001011011101,
       24'b001000010000010011011010,
       24'b000010100000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011011,
       24'b000001000000000011011000,
       24'b000000000000000011011001,
       24'b000000000000000011011011,
       24'b000011110000000011011001,
       24'b001100010001010011011100,
       24'b010111010100100011100010,
       24'b011111000110110011100101,
       24'b101001001001110111101011,
       24'b110111001101100111110011,
       24'b111111111111111111111001,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100001110111011110110,
       24'b010000100010011011011011,
       24'b000100010000100011010111,
       24'b100000110111001011100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b110111111101101011110100,
       24'b101011101010100011101110,
       24'b100011010111111111101000,
       24'b010110100100011011100000,
       24'b001011100001010011011011,
       24'b001001110000111011011011,
       24'b001111110010001011011011,
       24'b000010000000000011010110,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000011100000000011011001,
       24'b000010110000000011011001,
       24'b001000100000010011011011,
       24'b010010110011001111100001,
       24'b011100110110000111100110,
       24'b100101011000101011101001,
       24'b110001111100001111110001,
       24'b111101001111010111111000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111110011111100011111010,
       24'b110110111101100011110100,
       24'b101110001010111111101100,
       24'b111011101110110011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110011111100011111101,
       24'b010101100011111111011110,
       24'b000110100000111011011000,
       24'b010011010011000111100011,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b111011101110110111110101,
       24'b101110001011010011101101,
       24'b100010000111111011101001,
       24'b011101100110001111100011,
       24'b011011100101100111011101,
       24'b000111000000000011011001,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b000000000000000011011000,
       24'b001001010000001011010100,
       24'b001011000000110111011011,
       24'b000011000000000011011101,
       24'b001110110010001111011111,
       24'b011110000110011011100101,
       24'b101010011010001111101010,
       24'b101110011011010111101101,
       24'b111000101110001111110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b111000101110001111110010,
       24'b111011011110101011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b101111001011001111101010,
       24'b000011110000001011010010,
       24'b000000000000000011010010,
       24'b101010011001110111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100010000111011111100100,
       24'b001010100000111111010011,
       24'b010001000010011011011000,
       24'b111011011110101111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111000111110000111111000,
       24'b110000101011110011110011,
       24'b100110111000110111101010,
       24'b011001000101000111100011,
       24'b010011100011010111100000,
       24'b001100000001000111011110,
       24'b000011000000000011011000,
       24'b000000000000000011011011,
       24'b000000110000000011011001,
       24'b000000000000000011010111,
       24'b000000110000000011011001,
       24'b000011100000000011011001,
       24'b000111110000000011010111,
       24'b001111110010010011011100,
       24'b010110110100011111100010,
       24'b100001110111011111100111,
       24'b101101011010110011101110,
       24'b110111111101110011110110,
       24'b111111111111111111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100011100101011110010,
       24'b011101110111001111100000,
       24'b010011110011101111100000,
       24'b000111110000111111010110,
       24'b011011100101001011011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b110001111011111011110100,
       24'b000011110000000011011001,
       24'b000000000000000011011000,
       24'b011110000110000111100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111001011010011101101,
       24'b001000000001000011011000,
       24'b000111000000010011010111,
       24'b110011001100010011110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100011111001111111010,
       24'b110101111101001011110100,
       24'b101011111010011111101100,
       24'b100110111000111111011111,
       24'b011000100100111011011100,
       24'b001010000000110011011100,
       24'b000010110000000011011010,
       24'b000000000000000011010111,
       24'b000000000000000011011001,
       24'b000000000000000011011001,
       24'b000000000000000011010101,
       24'b000010000000000011010110,
       24'b000101000000000011011010,
       24'b001100110001010111100000,
       24'b010010100011011111100000,
       24'b100100000111111111100101,
       24'b110000001011011011101101,
       24'b110110111101100111110011,
       24'b111111011111111111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b110101001101010011110011,
       24'b110010011100001011110010,
       24'b110101101101011111110010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100001010010011101100,
       24'b000000000000000011010010,
       24'b000000000000000011011101,
       24'b000110000000000011011101,
       24'b000010110000000011011000,
       24'b110010001100000011110011,
       24'b111111111111111111111111,
       24'b111100011110111111111010,
       24'b001010100000100011011110,
       24'b000101110000100111011000,
       24'b011010010101010011011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011011100011111110101,
       24'b000101110000011011011101,
       24'b000001100000000011011000,
       24'b100110001000011111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111110111111010,
       24'b111101101111011111110110,
       24'b110000001011100011110000,
       24'b100000010111101011101010,
       24'b010110010100010011100001,
       24'b001011110001001111011100,
       24'b000111110000000011011011,
       24'b000001000000000011011001,
       24'b000010110000000011010110,
       24'b000101010000000011011010,
       24'b000101110000000011010110,
       24'b001011100001010111010101,
       24'b001001000000101011011010,
       24'b001010000000111111011010,
       24'b010111110100100011011111,
       24'b100001010111010011100100,
       24'b100111101001010111101000,
       24'b110010101100010011110000,
       24'b111100001110111111111001,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b101010001001101111101011,
       24'b001111100010111011011100,
       24'b000101000000000011011010,
       24'b000110000000000011011001,
       24'b000101110000000011011000,
       24'b001110010010111111011110,
       24'b110110001101000111110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101011111001111110111,
       24'b001110110001101111011100,
       24'b001000110000100011011110,
       24'b001010000000011011011111,
       24'b000000000000000011011011,
       24'b010100100011011011100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110000011111111100010,
       24'b000010100000001111011010,
       24'b010000110010010011011111,
       24'b111101101111010011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101001111001011111001,
       24'b001110110001100011011110,
       24'b000001100000001111011011,
       24'b011000100100100011100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111101,
       24'b111000111110001111110111,
       24'b101101011010111111101110,
       24'b100001010111100111100111,
       24'b011001000101000011100100,
       24'b001110110001111011011101,
       24'b001110110001101111011101,
       24'b000101000000000011011100,
       24'b000000000000000011010111,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b000010010000000011011010,
       24'b000101100000000011011011,
       24'b001101100001110111011101,
       24'b011100000110000111100101,
       24'b101100011010101011101011,
       24'b111000111110000011110000,
       24'b111001111110100011110101,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111111111110,
       24'b111111111111111111111110,
       24'b111101001111001011111011,
       24'b110001111100000111110001,
       24'b111100001110111011111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100011110111101011100111,
       24'b000000000000000011010100,
       24'b000001100000000011011100,
       24'b000000000000000011011011,
       24'b001111100010001011011110,
       24'b010110110011111011100100,
       24'b000000000000000011011000,
       24'b001011010000111011011000,
       24'b111100111111001011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110100100000011100101,
       24'b000100000000011011011011,
       24'b001010110000101111011111,
       24'b001000000000000011100000,
       24'b000100010000000011010111,
       24'b110011111100100111110001,
       24'b111111111111111111111111,
       24'b100010110111110111101000,
       24'b000000000000000011011001,
       24'b000010100000000011011011,
       24'b110011101100011111110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010111000100001011100011,
       24'b000000000000000011011001,
       24'b010000100010000111100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111010,
       24'b111000011110000111110101,
       24'b101110101011101111101110,
       24'b110100001100100111101011,
       24'b100101001000011111100111,
       24'b001111010010101111011110,
       24'b001001100000011011011011,
       24'b000010010000000011011000,
       24'b000000000000000011011001,
       24'b000000000000000011011001,
       24'b000000000000000011011001,
       24'b000000000000000011010111,
       24'b000000000000000011010111,
       24'b001000110000000011011010,
       24'b001111010010001111011111,
       24'b010111000100100011100010,
       24'b100011101000000111101000,
       24'b101111111011100111110000,
       24'b110111101101111011110101,
       24'b111111111111111111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111011111101,
       24'b011010010101000111100100,
       24'b000110100001000111011011,
       24'b000000000000000011010011,
       24'b101110101011000011101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101101011110110,
       24'b000011010000000011011000,
       24'b000100100000000011011101,
       24'b000101110000000011011101,
       24'b010110000100010011100000,
       24'b100001000111001011100011,
       24'b001110000001110011100000,
       24'b001000000000011011011111,
       24'b000000000000000011010111,
       24'b100000000110110111100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011111000110011111101010,
       24'b000000000000000011011011,
       24'b001010000000010011011101,
       24'b001010110000101011011111,
       24'b000011010000000111011101,
       24'b010101100011100011100001,
       24'b111111111111111111111111,
       24'b101111011011001111101111,
       24'b000011110000000011011000,
       24'b000000000000000011011010,
       24'b100101011000010011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100011111000000011101001,
       24'b000000000000000011011000,
       24'b001000000000001011011110,
       24'b111001011110001011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111110111111110011111000,
       24'b110101011101000111110100,
       24'b101010101010000011101101,
       24'b011101100110010011100100,
       24'b010001000010101111011101,
       24'b001000010000001011011010,
       24'b000001010000000011011000,
       24'b001010100000110011011010,
       24'b010000000010001111011100,
       24'b000001000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b000110000000000011011010,
       24'b010010110011001011100000,
       24'b010101100011110111100001,
       24'b011110000110101011100101,
       24'b101011101010011111101100,
       24'b111000001101111011110110,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b110001111100100111110000,
       24'b101000111001011111100101,
       24'b100001101000000111100110,
       24'b100110101001010111101011,
       24'b111010011110001011111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100110011101011100011,
       24'b000000000000000011010111,
       24'b000000000000000011011001,
       24'b100100000111111111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111101001000111101100,
       24'b000000000000000011011000,
       24'b000100110000000011011011,
       24'b010110000100010011100100,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b101001111001101111101100,
       24'b000000000000000011011100,
       24'b000101000000010011011011,
       24'b010010100010111011011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b101000111001011011101110,
       24'b000000000000000011011001,
       24'b001001110000001011011110,
       24'b001011100000111111011100,
       24'b000101010000000011011111,
       24'b000000100000000011011001,
       24'b110111111101100111110111,
       24'b111110011111100011110111,
       24'b001000110000000111010110,
       24'b000000100000000011011010,
       24'b011000010100100111100101,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100111010011111110000,
       24'b000000000000000011011001,
       24'b000000000000000011011001,
       24'b101101011010100111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101111111100111111001,
       24'b110011101100110011110001,
       24'b101010011010000011101101,
       24'b100000110111010111101000,
       24'b010101110100000011100000,
       24'b001110100001111011011110,
       24'b000101010000000011011011,
       24'b000000110000000011010110,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011010111,
       24'b001101110001110011011000,
       24'b011011110101011111100001,
       24'b011011010110010011101000,
       24'b100110111001000111101010,
       24'b110011111100101011110001,
       24'b111110001111101011111000,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000101101110111110110,
       24'b001111010011000011011101,
       24'b000001000000000011010111,
       24'b000001110000000011010101,
       24'b000100100000000011010101,
       24'b000010110000000011010100,
       24'b001000010000101011010111,
       24'b110101011100111111110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001011001011111101110,
       24'b000000000000000011010111,
       24'b000000000000000011011010,
       24'b010111010100001111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110001000100111101011,
       24'b000000000000000011011001,
       24'b000010100000000011011001,
       24'b100011010111101111101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101001111001111111010,
       24'b001000110000100011011011,
       24'b001101000000111111011011,
       24'b010000000010000011011100,
       24'b111000111101111011111010,
       24'b111111111111111111111111,
       24'b110110001101001111110101,
       24'b000110010000000011011011,
       24'b000010100000000011011101,
       24'b011010010100111111100011,
       24'b010111000100001111100000,
       24'b000000000000000011011000,
       24'b010011110010111011100010,
       24'b111111111111111111111010,
       24'b010010010010110111100000,
       24'b000000000000000011011010,
       24'b010001000010001111100001,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110111101010111110111,
       24'b000110010000000011011010,
       24'b000000000000000011011001,
       24'b011110000110001111100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111001101110001011110110,
       24'b101100101010100111101110,
       24'b100100001000001011101000,
       24'b011011010101100011100101,
       24'b010011010011100011011110,
       24'b000110110000000011011000,
       24'b000001100000000011010111,
       24'b000000100000000011011001,
       24'b000000000000000011011100,
       24'b000000000000000011011000,
       24'b000101100000000011010101,
       24'b000111010000000011011001,
       24'b000110110000000111011100,
       24'b010100010011011011100001,
       24'b011101010110001111100101,
       24'b100111001001001011101011,
       24'b110000101011101111101110,
       24'b111001001110001111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111110111111010,
       24'b110010111100100011110011,
       24'b101110001011011111110010,
       24'b110100111101001111110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101101111010111111010,
       24'b001110000001100111011010,
       24'b000000000000000011011001,
       24'b000110010000000011011111,
       24'b000001000000000011011001,
       24'b000001100000000011011010,
       24'b000101100000000011011110,
       24'b000111110000010011011010,
       24'b001111100010010011011011,
       24'b111100011110111011111011,
       24'b111111111111111111111111,
       24'b110100101100110011110011,
       24'b000101100000000011011011,
       24'b000100100000001011011101,
       24'b010001110010100111011111,
       24'b111111001111101011111110,
       24'b111111111111111111111111,
       24'b101101001010101011110000,
       24'b000001100000000011011000,
       24'b000011100000000011011100,
       24'b010101110011101111100000,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010011000010110111011111,
       24'b000101000000001111011011,
       24'b000100000000000011011000,
       24'b101101011010101011110001,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b001110110001100011100001,
       24'b000000000000000011011010,
       24'b011100000101010011101000,
       24'b101100101010011111101000,
       24'b000010000000000011011000,
       24'b000011100000000011010101,
       24'b111000111110000111110000,
       24'b100011000111101111101101,
       24'b000000000000000011011000,
       24'b001000110000001011011100,
       24'b111010011110010111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010010000010011111011110,
       24'b000010110000000111010110,
       24'b010110100100001111100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100010000111011111100100,
       24'b000000000000000011010001,
       24'b000111110000000011011000,
       24'b000000000000000011011001,
       24'b000000000000000011011011,
       24'b000000000000000011011011,
       24'b000001110000000011011001,
       24'b000110010000000011011001,
       24'b010101100100000011011110,
       24'b100000110111001111100011,
       24'b101010111010000011100101,
       24'b110000011011111011110011,
       24'b110111111110000011110111,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b100010010111110111101000,
       24'b001101010010001011011101,
       24'b000110110000000011011001,
       24'b000000110000000011011010,
       24'b000010110000000011011000,
       24'b010101110100100011100000,
       24'b111110001111011011111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100011010010111110000,
       24'b000000000000000011011000,
       24'b001001010000011111011110,
       24'b010000110010011011011011,
       24'b101011001010000111101101,
       24'b110001001011110011110010,
       24'b001101100001100111011111,
       24'b000111100000100011011110,
       24'b000000000000000011011000,
       24'b101001001001011011101111,
       24'b111111111111111111111111,
       24'b111100111111001011111010,
       24'b001011100000101111011111,
       24'b000100000000000011011101,
       24'b001001100000011111011011,
       24'b111001011110001111110111,
       24'b111111111111111111111111,
       24'b111010101110011111111001,
       24'b001001010000001011011101,
       24'b000011010000000011011110,
       24'b000110100000000011011100,
       24'b111001001110000011110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110010110010011101000,
       24'b000000000000000011011001,
       24'b000000010000000011011001,
       24'b100001000111000111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110100100000111100010,
       24'b000000100000000011011010,
       24'b001001110000100011011110,
       24'b111001011110001111110011,
       24'b010110100011111011100011,
       24'b000000000000000011011000,
       24'b011011000101001111100011,
       24'b101011111010010011101010,
       24'b000100100000000011011100,
       24'b000000100000000011011000,
       24'b101100111010100111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101000101111011100101,
       24'b001001110000101011010011,
       24'b010101000011101011011100,
       24'b111110001111011011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011111010010011110000,
       24'b000001000000000011011000,
       24'b001001100000100111011110,
       24'b001111000001111111100000,
       24'b010100100011110011100001,
       24'b011111110110111111100110,
       24'b101011111010100111101110,
       24'b110100011101000111110011,
       24'b111110111111101111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111011111101,
       24'b111110111111101011111011,
       24'b110111111101111011111001,
       24'b101111001011100111110001,
       24'b111010001110010111110110,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110000110000011100100,
       24'b000000000000000011010011,
       24'b000101010000000011011101,
       24'b000001100000000011011011,
       24'b000000000000000011011001,
       24'b000100100000000011011110,
       24'b000000000000000011010110,
       24'b011001010100110011100010,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b100101111000010111101110,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b011111000110100111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011011010000111101101,
       24'b000000000000000011010010,
       24'b000000000000000011010000,
       24'b011100110101111111100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011000010100101111100010,
       24'b000100010000000111011001,
       24'b000000000000000011011001,
       24'b101100001010011011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010001100010011111100001,
       24'b000011000000000011011101,
       24'b000010000000000011011010,
       24'b101101111010110111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101000111001011011101110,
       24'b000000010000000011011000,
       24'b000001110000000011011100,
       24'b010110010011111111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001100111010011100111,
       24'b000000000000000011010110,
       24'b000000010000000011011001,
       24'b111000111110001011111000,
       24'b110100101100101111110011,
       24'b000000000000000011011001,
       24'b000111000000000011011111,
       24'b011100100101111111100000,
       24'b010000000001110111011110,
       24'b000010010000100111011001,
       24'b100001100111010011101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110011000100111101001,
       24'b000100110000101111010111,
       24'b001011100001101111011001,
       24'b110100111100111011110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000001101110011110111,
       24'b001000010000000011011100,
       24'b000000000000000011011010,
       24'b100010110111101011101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111011111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111011101110110111110110,
       24'b111100001110111011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b100000110111000011100011,
       24'b001011000010000111010100,
       24'b000000000000000011010011,
       24'b101000101001010011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011011100011111110011,
       24'b000011000000000011011000,
       24'b001001110000011111011111,
       24'b000101100000000011011100,
       24'b011000010100100111100011,
       24'b011110100110010011100111,
       24'b001000110000000011011100,
       24'b000100100000000011011110,
       24'b000011000000000011010111,
       24'b110111011101100111110010,
       24'b111111111111111111111111,
       24'b100111011000110111101110,
       24'b000000010000000011011001,
       24'b000001010000010011011011,
       24'b011010010100111111100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010111110100111111000,
       24'b011110010110110111100100,
       24'b101001101010000111101100,
       24'b110111101101101011110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100100001000000011101000,
       24'b000111110000101011011001,
       24'b000011110000100111011001,
       24'b011101100110000011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011001110100111111100110,
       24'b000010000000000011011001,
       24'b000001010000000011011000,
       24'b100101001000010011101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010101100010011110010,
       24'b000011010000000011011010,
       24'b000001010000000011011110,
       24'b001101010001001111011111,
       24'b111111101111111111111011,
       24'b111111111111111111111111,
       24'b101110011010111111110000,
       24'b000010100000000011011010,
       24'b000000000000000011011001,
       24'b100111101000111111101110,
       24'b111111111111111111111110,
       24'b001101000001001111011101,
       24'b000000000000000011011100,
       24'b001100110001001011011110,
       24'b010011100011010011011110,
       24'b001001000001100111011010,
       24'b011000100100100111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111111011011011110000,
       24'b000010000000000011011000,
       24'b000000000000000011011000,
       24'b100110101000101011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111011111101,
       24'b001111010001111011011111,
       24'b000000000000000011011010,
       24'b010101100011101011100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111111111101,
       24'b101101011010101111101110,
       24'b011110010111000111100101,
       24'b011000100100111011100011,
       24'b000100010000101111010100,
       24'b100010010111011011101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001000111001011100111,
       24'b000110000000011011010011,
       24'b000110110000101011010110,
       24'b011110100110011111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100011110111111111101100,
       24'b000000000000000011011001,
       24'b000010100000001011011101,
       24'b010110110100011111100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100101011000011111101010,
       24'b000000000000000011010111,
       24'b000000000000000011010100,
       24'b011011100101100011100101,
       24'b111111111111111111111111,
       24'b101111101011010111110010,
       24'b000010100000000011011000,
       24'b001000110000100011011100,
       24'b001000000000110111011100,
       24'b111100111110111111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111011000110011101110,
       24'b000110000000101011011000,
       24'b001100010001110011011100,
       24'b011000010100100111100010,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b100110111000101111101100,
       24'b000000110000000011010110,
       24'b000000110000000011011011,
       24'b011001110101000111100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101011111010011111001,
       24'b010000010010001111011101,
       24'b000111000000101111011101,
       24'b000010110000000011011000,
       24'b110100111100110111110101,
       24'b111111111111111111111111,
       24'b110111111101101011110111,
       24'b000110110000000011011101,
       24'b000000000000000011011001,
       24'b010111010011111111100010,
       24'b111111111111111111111111,
       24'b101101011010100111110000,
       24'b000000000000000011010111,
       24'b001101000001000011011110,
       24'b001100110001000111011111,
       24'b000010100000000011011101,
       24'b001111010001100111011111,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100011111001111111010,
       24'b001010010000010011011100,
       24'b000000000000000011010111,
       24'b011100110101110111101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010110101010011100110,
       24'b000000000000000011011000,
       24'b001001110000010111011110,
       24'b111011101110110011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111001001110011011110110,
       24'b110100111100011111110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b001101000001011011011010,
       24'b000000000000000011010101,
       24'b000000110000000011011100,
       24'b000010010000000011010111,
       24'b100011010111110011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111101011010011110100,
       24'b000001100000000011011011,
       24'b000011100000000011011011,
       24'b001111110001111011011111,
       24'b111111101111111111111100,
       24'b111111111111111111111111,
       24'b100011110111111111101101,
       24'b000000000000000011011000,
       24'b000000000000000011011001,
       24'b100010010111001011101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101011111110101,
       24'b001011000001110111011010,
       24'b010101100101001111100000,
       24'b101010111001111011101101,
       24'b111111111111111111111111,
       24'b111110011111100011111100,
       24'b001011110000111011011101,
       24'b000011110000000011011011,
       24'b000010000000000011011011,
       24'b010000100011010011011110,
       24'b111110011111010111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101001100111011110011,
       24'b000011010000000011011001,
       24'b000011000000000011011101,
       24'b001101000000111111011110,
       24'b111110001111011111111010,
       24'b111111111111111111111111,
       24'b110010111100001111110100,
       24'b000011010000000011011100,
       24'b000011000000000011011101,
       24'b001110100001101011011101,
       24'b111110111111101111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010101000011100111100000,
       24'b010101010011100111011110,
       24'b011111110111001111011111,
       24'b101000111001011011101010,
       24'b111111111111111111111111,
       24'b111110111111101111111101,
       24'b010011100011001011100000,
       24'b000101100000110011011101,
       24'b001010110000111011011101,
       24'b111111011111110111111101,
       24'b111111111111111111111111,
       24'b001110110001101011100000,
       24'b000000110000000011011100,
       24'b000111110000000011011111,
       24'b000111100000000011100000,
       24'b000101000000000011011010,
       24'b110101101101000111110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010011000010111111100010,
       24'b000000000000000011011001,
       24'b010011100010111011100010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110011000101011101110,
       24'b000000000000000011011001,
       24'b000110100000000011011010,
       24'b110101101101000111110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b110110011101010111110011,
       24'b011001000101110011100000,
       24'b010010010010111111011111,
       24'b000111010000001111011011,
       24'b000010010000000011010110,
       24'b110111001101100011110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010111000100010011011111,
       24'b000100110000001111011001,
       24'b000111110000000011011111,
       24'b000101000000010011011100,
       24'b010101010011100011100000,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111001111110010111110111,
       24'b001000100000001011011110,
       24'b000100000000000011011110,
       24'b000101110000000011011011,
       24'b110111101101101011111000,
       24'b111111111111111111111111,
       24'b101100011010010111110000,
       24'b000001100000000011010111,
       24'b000101100000001011011100,
       24'b001111010010000111011111,
       24'b111111111111111111111011,
       24'b111111111111111111111111,
       24'b111111011111101111111100,
       24'b111111011111110011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001101001100111101011,
       24'b000000000000000011010110,
       24'b000110100000000011100001,
       24'b000000000000000011011100,
       24'b001100100010000011011101,
       24'b101111011011011111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111110111111101,
       24'b001100000000101111011111,
       24'b000011010000000011011101,
       24'b000101110000000011011010,
       24'b110001101011111111110100,
       24'b111111111111111111111111,
       24'b111011101110110011111010,
       24'b001001010000001011011101,
       24'b000100000000000011011101,
       24'b000110110000000011011101,
       24'b111000011101110111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100000101100111100111,
       24'b000011110000100011011100,
       24'b001110100011010111011100,
       24'b100000010110111111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100101101000100011100100,
       24'b001100010001011011011010,
       24'b000001100000000011011100,
       24'b110101001100111011110111,
       24'b111111111111111111111111,
       24'b101011101001111111101110,
       24'b000000000000000011010111,
       24'b001110110001100011011110,
       24'b001010100000101111011101,
       24'b000000100000000011011001,
       24'b101011011010001011101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101100110001011100101,
       24'b000000000000000011011010,
       24'b001000010000000011011100,
       24'b111001011110010011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111001011001011110011,
       24'b000010110000000011011010,
       24'b000101110000011011010100,
       24'b101100001010011111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110000111011101111110001,
       24'b000000000000000011010101,
       24'b000000100000000011011100,
       24'b000110100000000011011110,
       24'b000000000000000011011000,
       24'b100001100111001011101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b011101000101111011100001,
       24'b000100000000001011011000,
       24'b001001000000000111011111,
       24'b000101110000000011011111,
       24'b000111000000000011011001,
       24'b111000001101110111110110,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b010010010010110111011101,
       24'b000010010000000011011110,
       24'b000110100000011011011011,
       24'b110100001100101111110100,
       24'b111111111111111111111111,
       24'b111011101110110111111001,
       24'b000111100000000011011100,
       24'b000110000000000011100000,
       24'b000000100000000011011011,
       24'b011111010110111111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b011111000110011011100101,
       24'b000100000000000011010011,
       24'b001000010000000011011111,
       24'b000010000000000011011100,
       24'b000010100000000011010111,
       24'b011010100110001011100011,
       24'b111010101110001111111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110000110001011100011,
       24'b000001010000000011011001,
       24'b000000010000000011011000,
       24'b100110001000101011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010010010010101111100000,
       24'b000011000000000111011011,
       24'b000010010000000011011000,
       24'b101101011010110011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101010001001101111101101,
       24'b000001000000000011010111,
       24'b000000000000000011011001,
       24'b010101010011101011100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111111000111111101001,
       24'b000100010000011011010101,
       24'b001000000000110111010111,
       24'b101110111011001111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010000000001111011011111,
       24'b000111010000111111011010,
       24'b001101000001001111011101,
       24'b000000000000000011011001,
       24'b100001110111010111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001111001101011110000,
       24'b000000010000000011011010,
       24'b000001000000000011011001,
       24'b101101101010110011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010111110101011111000,
       24'b001001110000010011011100,
       24'b000000000000000011010111,
       24'b011100000101110011100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101001111010011111010,
       24'b001100000000101111011111,
       24'b000101000000000011011101,
       24'b001101000001100011011110,
       24'b000101010000000111011101,
       24'b001110010001011111011111,
       24'b111111011111111011111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110000110000111101000,
       24'b000010010000000011011010,
       24'b001001110000011011011111,
       24'b001010010000100011011111,
       24'b000010110000000011011000,
       24'b101101101010110011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101000101111111100110,
       24'b000000000000000011011011,
       24'b000101000000011111011001,
       24'b101000111001010111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110000110001011100101,
       24'b000000000000000011010110,
       24'b001000110000001011100000,
       24'b000000010000000011011001,
       24'b011100110110011111100011,
       24'b111110011111100011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b100110101000100111100100,
       24'b000010110000000011011000,
       24'b000000000000000011011100,
       24'b001010010000011011011111,
       24'b000000000000000011011010,
       24'b000111010000111111011010,
       24'b110001001011100011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100111010100011100111,
       24'b000111000000001011011000,
       24'b000000000000000011011001,
       24'b011110000110010011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110110110011111100111,
       24'b000000000000000011011000,
       24'b000000000000000011011000,
       24'b100000010110111011101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101111101001011110111,
       24'b001010010000101111011010,
       24'b000110110000100011011101,
       24'b001010010000011111011110,
       24'b111100011111000011111011,
       24'b111111111111111111111111,
       24'b110010011100000111110101,
       24'b000010110000000011011101,
       24'b000010010000010011010110,
       24'b100011111000000011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101011010100111101111,
       24'b000000000000000011011000,
       24'b001000000000000011011111,
       24'b000001100000000011011011,
       24'b010101010011101111100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101001100110011110111,
       24'b000100100000000011011011,
       24'b000000000000000011010111,
       24'b100110111000101111101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010100010011010111100011,
       24'b000000000000000011011000,
       24'b010001100010011111100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110100011111111100001,
       24'b000101000000000111011011,
       24'b001101100001011111011110,
       24'b001000000000000011100000,
       24'b000000000000000011010111,
       24'b101111101011010111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100000000110110011101101,
       24'b000001010000000011010111,
       24'b001001000000001011100000,
       24'b001010100000011111011110,
       24'b000000110000000011011010,
       24'b100100101000000111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111011000111011101111,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b010110010011111111100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111111011111001,
       24'b010000100010100011011010,
       24'b000000000000000011011010,
       24'b001000100000000011100000,
       24'b000000000000000011011001,
       24'b001111010010010011011011,
       24'b101011111010100011101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010101100001111110001,
       24'b010011000011111111100000,
       24'b000000000000000011010111,
       24'b000110110000000011011111,
       24'b000101000000000011011100,
       24'b000000000000000011010111,
       24'b110001011011100111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101101010110011110001,
       24'b001101010001011111011000,
       24'b000101110000101011011100,
       24'b010001110010101111100010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b101100111010100011101111,
       24'b000000110000000011011001,
       24'b000000110000000011011011,
       24'b010101110011101111100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010001100010011011100000,
       24'b000011000000001111011100,
       24'b000010010000000011011000,
       24'b110001001011101111110010,
       24'b111111111111111111111111,
       24'b111100011111000111111001,
       24'b001011000000100011011100,
       24'b000000000000000011011011,
       24'b010011110011001011100010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010000010010000011011111,
       24'b000001110000000011011101,
       24'b000100010000000011011110,
       24'b000101000000000011011011,
       24'b111010111110101011111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100111111001111111010,
       24'b001001110000000111011110,
       24'b000000000000000011011000,
       24'b011011010101011011100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110000110010011101000,
       24'b000001010000000111011000,
       24'b001010110000010011011110,
       24'b111011001110101011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100010110111101011101010,
       24'b000000110000001011011001,
       24'b001001010000000011011110,
       24'b001000010000000011100000,
       24'b000001110000001011011001,
       24'b011011000101001011100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100011110111111011101100,
       24'b000000000000000011011000,
       24'b001110100001110011011010,
       24'b001011000000101111011100,
       24'b000001000000000011011011,
       24'b011000010100100111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111111011100011110001,
       24'b000101010000001111011001,
       24'b000100010000001011011101,
       24'b001110100001011011100000,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011101110101111111010,
       24'b010001100011011111011111,
       24'b000000000000000011010110,
       24'b000101100000000011011101,
       24'b000100010000000011011011,
       24'b000000000000000011011000,
       24'b011000110101100011100010,
       24'b111110001111010111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b100110101001001011101010,
       24'b000011110000000011011010,
       24'b000011100000000011011101,
       24'b000001000000000011011101,
       24'b001000010000010111011010,
       24'b111100011110111011111001,
       24'b111111111111111111111111,
       24'b110111101101101011111000,
       24'b001011000000111011011100,
       24'b010010010010011011011100,
       24'b001000110000001111011010,
       24'b111001101110001111110101,
       24'b111111111111111111111111,
       24'b110110101101011111110110,
       24'b000101100000000011011011,
       24'b000011000000000011011100,
       24'b001010010000110111011101,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010011100011001111100010,
       24'b000011000000000011011101,
       24'b000011100000000011010111,
       24'b101110001010111011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010011010011000011100000,
       24'b000000000000000011011011,
       24'b001010110000101011011111,
       24'b111110001111100011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101011010101011110000,
       24'b000000000000000011010010,
       24'b000011010000000011011000,
       24'b001001110000111111011011,
       24'b110101001100111111110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b011001000100110011100001,
       24'b000010000000000111011001,
       24'b001110010001110011011110,
       24'b111110011111100111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111001000110111101011,
       24'b000010100000001011010111,
       24'b000010110000000011011001,
       24'b101100101010100011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100001010001111110001,
       24'b000000010000000011011010,
       24'b001010010000001111011110,
       24'b001001100000010011011111,
       24'b000111110000000011011110,
       24'b000110000000000011011011,
       24'b111010011110011111111000,
       24'b111111111111111111111111,
       24'b100110111000100111101110,
       24'b000000000000000011011001,
       24'b010111000100010011100000,
       24'b010010000010101111100000,
       24'b000001010000000011011101,
       24'b001110000001010111011111,
       24'b111110101111100111111011,
       24'b111111111111111111111111,
       24'b111011111110110111111000,
       24'b001100010000110111011011,
       24'b000110100000001111011100,
       24'b000110110000000011011011,
       24'b110111101101101011110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b100010011000000011100111,
       24'b001000010000111111011001,
       24'b000000110000000011011001,
       24'b000111010000000011100000,
       24'b000000000000000011011001,
       24'b001101110010001011011001,
       24'b111011001110101111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011101100010111110001,
       24'b001001110001101011011011,
       24'b001011010000110111011110,
       24'b000000000000000011011000,
       24'b100010100111100111101000,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b001110000001011111100000,
       24'b001001110000110111011111,
       24'b000110010000000011010111,
       24'b101010011001110011101110,
       24'b111111111111111111111111,
       24'b111110101111110011111011,
       24'b001101100001000111011101,
       24'b000011010000000011011101,
       24'b000101100000011011011101,
       24'b100000010111000111100111,
       24'b110111001101011111110001,
       24'b101001011001100011101101,
       24'b000110100000001111011110,
       24'b000110100000000011011111,
       24'b001001110000011011011001,
       24'b111000011101111011110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101100110001011101000,
       24'b000000000000000011010100,
       24'b000000000000000011010001,
       24'b101110111011001011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111010,
       24'b101000001001001011101000,
       24'b110001101100000011110001,
       24'b111101001111010111111001,
       24'b111111001111101011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111111001001011100111,
       24'b000000110000000011010110,
       24'b001001010000010111011011,
       24'b111000111110000011110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110001101001011110110,
       24'b000111110000010111011000,
       24'b000000100000000011011010,
       24'b100011000111110111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000111101110111110111,
       24'b001001110000110111011011,
       24'b000101010000001111011111,
       24'b001111110010000111011100,
       24'b001011000000101011011101,
       24'b000001110000000011011000,
       24'b101000001001001011101011,
       24'b111111111111111111111111,
       24'b101001011001100011101111,
       24'b000000000000000011011000,
       24'b011000000100011111100011,
       24'b011000000100011011100010,
       24'b000010000000000011011101,
       24'b000110010000000011011100,
       24'b110110111101011111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010100110011011111100100,
       24'b000100100000000111011010,
       24'b000010010000000011011000,
       24'b101010001001101011101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010111110100111110101,
       24'b010110110100100011100000,
       24'b000000000000000011010111,
       24'b000110010000000011100001,
       24'b000000000000000011011000,
       24'b010110000011101111011100,
       24'b111111101111111011111100,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b111101011111001111111010,
       24'b101111101011101111101111,
       24'b110110111101011011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001111001011111101101,
       24'b000011100000100111011000,
       24'b000001100000000011011011,
       24'b010010110010111111011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b011001000100110111100011,
       24'b000000000000000011011011,
       24'b001100000001010011011010,
       24'b110010011100001011101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100100011000001011100111,
       24'b000000000000000011010111,
       24'b001010100000011011100001,
       24'b000011110000000011011011,
       24'b001000010000000011010111,
       24'b000011010000000011011010,
       24'b000111100000000011100000,
       24'b000000000000000011011000,
       24'b010111010100010011100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100111010100011110000,
       24'b010101100100100111011110,
       24'b100101011000101011100100,
       24'b110110001101000111110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111101011010111110000,
       24'b000011000000000011011010,
       24'b001000000000011111011010,
       24'b110101011101000011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111101111111101,
       24'b010000000001111111011110,
       24'b000010100000000011011000,
       24'b011010010101000011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b010001000010010111011110,
       24'b000001000000000011011100,
       24'b010111100100011011100001,
       24'b010110000011111111011111,
       24'b000111100000110011011000,
       24'b010100100011001111011100,
       24'b111111111111111111111111,
       24'b101110011011000011110010,
       24'b000000000000000011010111,
       24'b011010000101000011100100,
       24'b011111010110100111100011,
       24'b000001010000000011011100,
       24'b000001000000000011011000,
       24'b101100111010011111101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110000110001111101001,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b011111010110100111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001100111100111100111,
       24'b000110100000001111010111,
       24'b001011110000110111011110,
       24'b000001000000000011010100,
       24'b101001011001100011101101,
       24'b111111111111111111111111,
       24'b101100111010011111101110,
       24'b000110010001001011010111,
       24'b000000000000000011010001,
       24'b100011100111111011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011001110100111110111,
       24'b001011110001011111011000,
       24'b000010010000000011011100,
       24'b001100100000111111100000,
       24'b111110011111101011111100,
       24'b111111111111111111111111,
       24'b100110001000100111101100,
       24'b000000000000000011010111,
       24'b000110110000111011011100,
       24'b100101001000011011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111110111111100,
       24'b010100000011101011011111,
       24'b000000000000000011010100,
       24'b000000000000000011011010,
       24'b000000000000000011011101,
       24'b000000000000000011011001,
       24'b000000000000000011010111,
       24'b010000100011010111011111,
       24'b111010111110100011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111001001110000111110110,
       24'b001010100000010111011011,
       24'b000000010000000111011001,
       24'b100001000111000111101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010111100100011011100010,
       24'b000000000000000011011000,
       24'b001110110001100011100001,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010110101010011100110,
       24'b000000000000000011011001,
       24'b010110100011110011100101,
       24'b100011100111110111101001,
       24'b000101110000001011011010,
       24'b000010110000000011011001,
       24'b111011011110101111111000,
       24'b110110111101011011110111,
       24'b000000100000000011011001,
       24'b011000110100101111100110,
       24'b101001011001011111101101,
       24'b000110010000001011011011,
       24'b000000100000000011011010,
       24'b011111110110101011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111011000111011101100,
       24'b000000000000000011011000,
       24'b000000000000000011011011,
       24'b010101110011110011100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110011111100111111001,
       24'b111100111111001011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101100110000011100010,
       24'b000101100000010011011010,
       24'b000010100000000011011011,
       24'b010110010011111111100011,
       24'b111111111111111111111111,
       24'b110010111100010011110001,
       24'b000000000000000011011000,
       24'b000000100000000011011101,
       24'b010100110011110111011101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111001101011011110001,
       24'b000110110000100011011000,
       24'b000100010000000011011110,
       24'b001100100001001011011111,
       24'b111110001111100011111011,
       24'b111111111111111111111111,
       24'b110000111011110011110101,
       24'b000110000000000111011010,
       24'b000010100000000011011100,
       24'b000110000000000011011110,
       24'b111101111111011011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b100100011000110011101000,
       24'b010100000100001011100000,
       24'b010100010011101111011111,
       24'b011010100101110111100011,
       24'b101011011010101111101101,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111110111111100,
       24'b010011010011000111011110,
       24'b000000000000000011010111,
       24'b010011100011000111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011111000110100111101000,
       24'b000001110000000011011001,
       24'b001011110001001011011001,
       24'b110101001100110111110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100011100111110111101010,
       24'b000000000000000011011000,
       24'b000111110000000011011111,
       24'b101100101010011111101011,
       24'b010100010011010011100001,
       24'b000000000000000011011011,
       24'b100100101000000011101010,
       24'b111001001110000111110101,
       24'b000000000000000011011010,
       24'b010011010011001011100100,
       24'b110010001011111011110100,
       24'b001010010000001111011111,
       24'b000011000000000011011010,
       24'b010101000011100011100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111000111110000011110011,
       24'b001001010001000011011000,
       24'b001000010001010011011110,
       24'b010011100011000111100000,
       24'b111100111111001011111011,
       24'b111111111111111111111111,
       24'b110100001100100011110011,
       24'b011000000101110011100001,
       24'b001000010001101011011000,
       24'b100111011001000011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101001100110111110100,
       24'b000100100000000011011011,
       24'b000010110000000011011110,
       24'b001110010001101111011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b001100110000111011011111,
       24'b000011010000000011011100,
       24'b000110110000000011011011,
       24'b011111000110011111100110,
       24'b101000001001001111101010,
       24'b010000110010101011011111,
       24'b000101010000000011011101,
       24'b000000000000000011011001,
       24'b010100000011010111100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111001101110001111111000,
       24'b000011110000000011011000,
       24'b000000000000000011010100,
       24'b000111110000000011010100,
       24'b110111111101101111110101,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b110101111101010011110100,
       24'b111010101110100011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101100110001011100111,
       24'b000000000000000011010111,
       24'b001010010000011011011111,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101111010111011110001,
       24'b000010010000000011011001,
       24'b000001110000010011011000,
       24'b101010001001101111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101101010111011110001,
       24'b000000000000000011010111,
       24'b000000010000000011011010,
       24'b101111001011001111110000,
       24'b100100011000000011101011,
       24'b000000000000000011010111,
       24'b010010000010010011100001,
       24'b101111101011011111110010,
       24'b000101100000000011011110,
       24'b001101000001000111011111,
       24'b110111101101101111110100,
       24'b001111110010000011100010,
       24'b000010000000000011011101,
       24'b001100110001001011011100,
       24'b111011111110111111111000,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b010000100010001111011110,
       24'b001101000001110011011101,
       24'b010001010010110111011010,
       24'b110001111011111111110011,
       24'b111111111111111111111111,
       24'b101100001010010111101111,
       24'b000000000000000011010100,
       24'b000100100000000011011000,
       24'b100011000111101111100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111111111111001,
       24'b001000100000000011011011,
       24'b000110000000100111011011,
       24'b001100110001001111011110,
       24'b111101101111010111111100,
       24'b111111111111111111111111,
       24'b101000011001001111101100,
       24'b000000000000000011010110,
       24'b000110110000000011011110,
       24'b000001100000000011011001,
       24'b000000100000000011011001,
       24'b000100100000000011011110,
       24'b000010000000000011011110,
       24'b000000000000000011010100,
       24'b110001101011111011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111101111111100,
       24'b100101011000011011101001,
       24'b101000111001100111101001,
       24'b111000011101111011110010,
       24'b111110011111100111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110001111011011111001,
       24'b111010001110010111110101,
       24'b101111111011011111101111,
       24'b100110111001000111101011,
       24'b011011110101110011100100,
       24'b001111010010001111011101,
       24'b000000000000000011010100,
       24'b011100100101111111100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110001000100111101111,
       24'b000010010000000011011001,
       24'b001100100001000011011010,
       24'b110011101100011111110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011011110101111111000,
       24'b001001010000001111011110,
       24'b000000000000000011011000,
       24'b100001100111010011101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100001110111111110111,
       24'b001111000001111011011100,
       24'b000000000000000011011001,
       24'b100011100111110111101100,
       24'b111000111101111111110110,
       24'b000100100000000011011100,
       24'b000100000000000011011110,
       24'b011110000110001011100010,
       24'b001110000001001011011111,
       24'b000100110000000011011101,
       24'b111101101111100011110111,
       24'b011011110101100011100111,
       24'b000011110000010011011010,
       24'b001000000000011111011000,
       24'b110010111100010011110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010101010011100011100100,
       24'b000000000000000011011010,
       24'b000000000000000011010101,
       24'b101001101001100111101101,
       24'b111111111111111111111111,
       24'b111100011110111111111010,
       24'b000111000000000011011100,
       24'b000111110000011011011100,
       24'b001000110000111111011100,
       24'b101011111010011011101110,
       24'b111000001101110011110111,
       24'b011101100110000111100110,
       24'b000101010000001011011100,
       24'b000110010000101111011001,
       24'b010001000010100011011110,
       24'b111111001111101111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b011111110110100111100101,
       24'b000000110000000011010111,
       24'b000000000000000011011000,
       24'b000000010000000011011001,
       24'b000010010000000011011010,
       24'b001011010010000011011100,
       24'b101110011010101011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b111101101111011111111010,
       24'b110011001100100011110011,
       24'b100100111000110011100111,
       24'b111011001110100111110111,
       24'b111100011110111011111001,
       24'b001001110000100011010111,
       24'b000001000000000011011001,
       24'b000000000000000011011000,
       24'b000000000000000011010100,
       24'b000000000000000011010111,
       24'b000000000000000011010111,
       24'b010111100100011011011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111011011010011110011,
       24'b000100100000000011011011,
       24'b001000010001001111010110,
       24'b100101111000100011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010001100010010011100001,
       24'b000000000000000011011000,
       24'b010100010011011011100001,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b011000100100101011011111,
       24'b000000000000000011011001,
       24'b010001110010011111100011,
       24'b111111111111111111111101,
       24'b010100100010111111100001,
       24'b000000000000000011011100,
       24'b001101010001010111011100,
       24'b010000010010010111011100,
       24'b001100110001101011011110,
       24'b111110111111101111111101,
       24'b101001101001011111101111,
       24'b000000100000000111011001,
       24'b000000100000000111011000,
       24'b100110111000110011101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100000100111000111100111,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b011111110110101111101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110100110000111100101,
       24'b000000000000000011010111,
       24'b000101110000000011011110,
       24'b000101100000000011011011,
       24'b001001000000000011011100,
       24'b000100100000000011011011,
       24'b000110100000000011100001,
       24'b000000000000000011010101,
       24'b100110011000110011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100011100111011110100,
       24'b100110111001010111101010,
       24'b100111111001011011101001,
       24'b110000111100001011110001,
       24'b111111101111110011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101011111010111111100,
       24'b111000001101110011110011,
       24'b101011101010011111101101,
       24'b100001000111001111100100,
       24'b010111100100011111011111,
       24'b001100010001010011011110,
       24'b000000110000000011011000,
       24'b000000000000000011001011,
       24'b100011010111110011100111,
       24'b111111111111111111111111,
       24'b001101010001001011100001,
       24'b000001010000000011011100,
       24'b001110110010001011011111,
       24'b011101110110011111100110,
       24'b101010001001111111101101,
       24'b110100101100111011110101,
       24'b111011101110101011110111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100011111000011111000,
       24'b001001100000010011011100,
       24'b000000000000000011011001,
       24'b011110000110011111100001,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010010101000111100100,
       24'b000000000000000011011000,
       24'b001010000000011011011110,
       24'b111100001111000011111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011011100101100011100101,
       24'b000110100000111011011001,
       24'b001000010000000011011010,
       24'b111111111111111111111010,
       24'b101100111010100011101110,
       24'b000000000000000011011000,
       24'b000111100000000011011111,
       24'b001010000000101011011110,
       24'b001100000001011111011010,
       24'b111100001110111111111100,
       24'b110100011100101111110100,
       24'b000000100000000011011000,
       24'b000000000000000011011011,
       24'b011010010101001011100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101101010110111110000,
       24'b000001110000000011010111,
       24'b000001110000000011011100,
       24'b010011000010110111100001,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111100101111000111111010,
       24'b001110100010011011011100,
       24'b000000000000000011010111,
       24'b000000000000000011011011,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011010110,
       24'b011011000101011111100010,
       24'b111111111111111111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000001101110011110110,
       24'b110000111011110111110011,
       24'b100001010111110111100111,
       24'b110010001011111111110010,
       24'b111100101111000011111010,
       24'b000111110000000011011001,
       24'b000000000000000011010101,
       24'b000000000000000011010101,
       24'b000001110000000011011011,
       24'b001010100000011011011101,
       24'b001101010001011011011110,
       24'b001011100010001011011011,
       24'b100111011001000111100101,
       24'b111111111111111111111111,
       24'b011011100101011011101001,
       24'b000000000000000011010101,
       24'b011001110101001011100000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010101100011100111100011,
       24'b000000000000000011011001,
       24'b010011000010110011011110,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111111001000111101110,
       24'b000000000000000011011000,
       24'b000101000000000011011011,
       24'b110100011100101111110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001011001100011101101,
       24'b000100010000100111011001,
       24'b000001110000000011011000,
       24'b110011011100011111110100,
       24'b111111111111111111111111,
       24'b000111010000000011011100,
       24'b000110000000000011011110,
       24'b000110110000000011011111,
       24'b000011110000000011010111,
       24'b111001101110010111110110,
       24'b111101111111011111111011,
       24'b000110010000000011011001,
       24'b000000110000000011011101,
       24'b010001010010011111100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111010101110100111110111,
       24'b001001010000010111011011,
       24'b000010110000000011011100,
       24'b000101110000000011011101,
       24'b111001001110001011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111011111111010,
       24'b011111110111100111101000,
       24'b010101110100011111100010,
       24'b010110110100100111100010,
       24'b011101100110110011100111,
       24'b101111101011010011101111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111101111111011111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101001111001111111001,
       24'b100111111001000011101011,
       24'b011110100110101011100110,
       24'b100001110111010111100110,
       24'b001011110001001111011101,
       24'b000000000000000011011001,
       24'b000000000000000011010000,
       24'b010000000010001011011101,
       24'b111111111111111111111010,
       24'b001111010001111111011101,
       24'b010000010010100011011111,
       24'b010011100011001111100100,
       24'b000100010000000011011111,
       24'b000101110000100111011010,
       24'b101110011011000111101100,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b100011010111110111101001,
       24'b000000000000000011010111,
       24'b001100000000110111011110,
       24'b111100101111001011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011110110110011111100111,
       24'b000000000000000011011000,
       24'b001000000000000011011101,
       24'b111001111110011011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011111100011111110110,
       24'b000011010000000011011010,
       24'b000000100000000011011000,
       24'b101001011001011111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100001100100011110100,
       24'b000010100000000011011001,
       24'b000001010000001111011000,
       24'b100101011000010111101100,
       24'b111111111111111111111111,
       24'b011101000101110011100011,
       24'b000000000000000011011011,
       24'b001000110000000111100000,
       24'b000101100000000111011000,
       24'b110010011100001111110101,
       24'b111111111111111111111111,
       24'b001111100001101111100000,
       24'b000001100000000011011011,
       24'b001001110000001111011101,
       24'b111010011110011011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b001010110000100011011100,
       24'b000000000000000011010101,
       24'b000011000000000011010111,
       24'b110010001100001111110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111101111111001,
       24'b111101101111011011111010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101011111010111111010,
       24'b000101000000000011011000,
       24'b000000000000000011011000,
       24'b000101100000000011011010,
       24'b000110000000000011010110,
       24'b000111100000001011011001,
       24'b010000110011011011011111,
       24'b100100011000000111101001,
       24'b111111101111111111111100,
       24'b111001011110001111110110,
       24'b111111111111111111111101,
       24'b111110101111101011111010,
       24'b001011110001001011011100,
       24'b000000000000000011010111,
       24'b101110001011000011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010101100001011110000,
       24'b000011100000000111011011,
       24'b000000010000000011011001,
       24'b110001001011110011110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101000101001010011101100,
       24'b000000000000000011010111,
       24'b000000110000000011011001,
       24'b101100101010100111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011101110110111111001,
       24'b001010100000010011011101,
       24'b000000000000000011011001,
       24'b011011000101010111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110111111101111111010,
       24'b001100010000110111011111,
       24'b000011100000011011011000,
       24'b011001100100111011100010,
       24'b111111111111111111111111,
       24'b110011111100101011110010,
       24'b000010100000000011011000,
       24'b001001010000001111011111,
       24'b000001110000000011011011,
       24'b101100011010011011110001,
       24'b111111111111111111111111,
       24'b010101110011110111100110,
       24'b000000000000000011010100,
       24'b000000000000000011010010,
       24'b101010111001111111101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101100001010010111101111,
       24'b101001001010001111101110,
       24'b110110111101101011110101,
       24'b111110001111011111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110001111100011111100,
       24'b100100000111111011100111,
       24'b001010010001111011010111,
       24'b100011111000000111101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011001110100111011100101,
       24'b000000000000000011011001,
       24'b001110100001110111100000,
       24'b101111111011100111101111,
       24'b111010001110011011110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111101111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010100010011010011100000,
       24'b000000110000000011010111,
       24'b100001010111010011100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110101111101011111011,
       24'b010000100010001011011101,
       24'b000010010000001111010110,
       24'b100011010111110111101010,
       24'b111011001110101111110111,
       24'b100111111001100111101010,
       24'b100011010111100111100110,
       24'b111110111111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110011101001011110111,
       24'b000110000000000011011010,
       24'b000000000000000011011010,
       24'b100001000111000111101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010101100011101011100001,
       24'b000001010000000011011010,
       24'b001110000001011111011111,
       24'b111111101111110111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b011100100101110111100011,
       24'b000000000000000011011011,
       24'b001011000000011011011110,
       24'b111111001111110011111101,
       24'b111111111111111111111111,
       24'b001111100001111011011100,
       24'b000000000000000011010111,
       24'b000000000000000011010000,
       24'b100100111000010011100111,
       24'b111111111111111111111111,
       24'b101001011001011111101100,
       24'b011000110101111111100001,
       24'b101001101010010011101101,
       24'b111000111110000011110111,
       24'b111111111111111011111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111011111101,
       24'b111111111111111111111101,
       24'b111011101110110011111000,
       24'b110000111100000011110011,
       24'b100111011001001111101011,
       24'b011110100110101111100101,
       24'b100000111000000011100110,
       24'b111011001110010111110110,
       24'b111111111111111111111111,
       24'b111111011111110111111110,
       24'b001010100000100011011010,
       24'b000000000000000011010100,
       24'b011000000100100011100011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110001000100011101101,
       24'b000000000000000011010111,
       24'b010000010001110111100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011011110101100011100110,
       24'b000000000000000011010110,
       24'b010010000010101011011101,
       24'b111111101111111011111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010011110011001011100001,
       24'b000011000000000111011100,
       24'b001011110000110111011111,
       24'b001010100000011011011011,
       24'b000000000000000011010101,
       24'b000000000000000011010001,
       24'b110011101100100011110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b001110100001010111100000,
       24'b000000000000000011011000,
       24'b011010100101000111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001100111001111101001,
       24'b000000000000000011011001,
       24'b000111000000000011011100,
       24'b111000011101110011110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001000111001111100111,
       24'b000000000000000011010010,
       24'b000000000000000011010100,
       24'b110010011100001011110011,
       24'b111111111111111111111111,
       24'b101010011001110011101101,
       24'b010110010101100011100000,
       24'b100101001000111111101000,
       24'b110111101101101111110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100011111000011111001,
       24'b111000101101111011110100,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b011100010101101011100000,
       24'b000110100000110011011000,
       24'b001000010000000111011011,
       24'b000000000000000011010110,
       24'b000000000000000011010110,
       24'b000000000000000011011000,
       24'b001000110000110111011010,
       24'b111001011110000111110110,
       24'b111111111111111111111111,
       24'b100001000111000011101001,
       24'b000000000000000011010111,
       24'b010000100010001011011111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110011011000111110010,
       24'b000000010000000011011000,
       24'b000011010000000011011010,
       24'b110011101100100011110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101010101001101111101110,
       24'b000000000000000011011000,
       24'b001001010000011111011010,
       24'b111001011110001011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100010101101011100101,
       24'b000000000000000011011010,
       24'b000110100000000011011111,
       24'b000100010000000011011011,
       24'b010000100010011111011111,
       24'b010110000101000011100000,
       24'b110100011100100111110011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110010011111011100011,
       24'b000000000000000011010111,
       24'b010000010001111111100000,
       24'b111111001111101111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101010011001110111110000,
       24'b000000000000000011011000,
       24'b000001110000000011011001,
       24'b101110101011000111110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110111011000111110000,
       24'b010101000100111011011111,
       24'b100100001000101111101000,
       24'b111000111101111111110101,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b101101011010101011101111,
       24'b010011110100100111100000,
       24'b001000000000111111011001,
       24'b010000110010010111011001,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b010110110100000111100010,
       24'b000000000000000011011000,
       24'b001011010000110011011110,
       24'b010110010011110111100011,
       24'b011010010101010011100010,
       24'b001001010000000011011101,
       24'b000000000000000011011001,
       24'b011010000101000011100011,
       24'b111111111111111111111111,
       24'b101011101010001011110000,
       24'b000000000000000011011000,
       24'b001000100000000111011011,
       24'b111010101110101011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111001111110010011110111,
       24'b001000110000010011011010,
       24'b000000000000000011010111,
       24'b101001011001011111101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111110011111000,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100111100110111110101,
       24'b000100010000000011011100,
       24'b000001000000000011011011,
       24'b110000101011100111110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001001001011011101101,
       24'b000000000000000011011000,
       24'b000110010000000111011100,
       24'b101101111011000111101110,
       24'b111111101111111111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001100111010011101000,
       24'b000000010000000011011010,
       24'b000110110000000111011001,
       24'b110011101100011011110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100011100101111110010,
       24'b000100100000000011011010,
       24'b000000000000000011011000,
       24'b100001110111010111101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111100101111001011110111,
       24'b110000101011110111101110,
       24'b100100111000100011101001,
       24'b011000110101100111100011,
       24'b111001011110000011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100010101101111101000,
       24'b000000000000000011010100,
       24'b000100010000000011011100,
       24'b000101000000000011011011,
       24'b110101111101000111110110,
       24'b111111111111111111111111,
       24'b100111011000111011101110,
       24'b000000000000000011011000,
       24'b001000010000000011011101,
       24'b111110101111101011111010,
       24'b111111111111111111111111,
       24'b100000010110110111100111,
       24'b000000000000000011010111,
       24'b001100100000110011011111,
       24'b111111111111111111111111,
       24'b111000101101111111110111,
       24'b000011010000000011011001,
       24'b000001110000000011011000,
       24'b101111001011001111101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010011000010111011100001,
       24'b000000110000000011011010,
       24'b010101010011101111100011,
       24'b100011100111111011101010,
       24'b011001110101001011100001,
       24'b010011110011011011011010,
       24'b111000001101101111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100111111001111111010,
       24'b001011100000100111011101,
       24'b000000000000000011011000,
       24'b100100000111111011101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011111100100111110110,
       24'b000100100000000011011011,
       24'b000001000000000011011001,
       24'b110011101100011011110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111001011001111110001,
       24'b000001110000000011011011,
       24'b000000100000000111011000,
       24'b101010101001110011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111110011111010,
       24'b001110110001011011100000,
       24'b000000000000000011011001,
       24'b010101100011101111100010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111111111011,
       24'b110110101101100011110111,
       24'b110110011101010111110101,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101001100111111110001,
       24'b000001100000000011010101,
       24'b000000000000000011011001,
       24'b000000000000000011010110,
       24'b100011000111101011101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100101101000010011101111,
       24'b000000000000000011011010,
       24'b001010100000100011011110,
       24'b000010010000000011011000,
       24'b101011001001111011110001,
       24'b111111111111111111111111,
       24'b110011011100011111110101,
       24'b000011100000000011011001,
       24'b000010100000000011011010,
       24'b110100011100101011110101,
       24'b111111111111111111111111,
       24'b101111111011011011110010,
       24'b000000000000000011011000,
       24'b000100010000000011011011,
       24'b111010011110011011111001,
       24'b111111111111111111111111,
       24'b001111000001100011011111,
       24'b000000000000000011011000,
       24'b011110100110010111101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100010101110011101001,
       24'b000000100000000011011011,
       24'b000110110000000011011110,
       24'b000000000000000011010111,
       24'b000000000000000011010101,
       24'b000000000000000011001111,
       24'b101100001010010011101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010111000100001111100000,
       24'b000000000000000011010111,
       24'b010110010011111111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011111110111011111001,
       24'b001100000000111011011101,
       24'b000000000000000011010111,
       24'b100100000111111111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111000101110000011111000,
       24'b000111100000000011011011,
       24'b000000000000000011011000,
       24'b100000010110111111101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011011010101011111100110,
       24'b000000000000000011010111,
       24'b001110100001011111011111,
       24'b111111101111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111101000111011101000,
       24'b001100110001111111011011,
       24'b000101010000000011011101,
       24'b000101000000000011011010,
       24'b010000110011011111011110,
       24'b111001101110001011110110,
       24'b111111111111111111111111,
       24'b111110011111100011111101,
       24'b001100100001000111100000,
       24'b000101110000001011011100,
       24'b000101000000001111011111,
       24'b001100110001001011011110,
       24'b111111001111110111111100,
       24'b111111111111111111111111,
       24'b101001001001011011101110,
       24'b000000110000000011011000,
       24'b001000110000000011011111,
       24'b000000000000000011011001,
       24'b100001100111001011101010,
       24'b111111111111111111111111,
       24'b111100011111000011111000,
       24'b001011000000011111011100,
       24'b000000000000000011010111,
       24'b100110101000101011101100,
       24'b111111111111111111111111,
       24'b111000101101111011110110,
       24'b001011010001010111011011,
       24'b000000000000000011010111,
       24'b101000011001001011101101,
       24'b111111111111111111111111,
       24'b011001010100110011100110,
       24'b000000000000000011010110,
       24'b010100110011011111100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100101101000100011101011,
       24'b000000000000000011011001,
       24'b001000100000001011011110,
       24'b011000010100101111100011,
       24'b100000000110111111101001,
       24'b101001111010001011101101,
       24'b111001101110001011110111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100001000111001011101011,
       24'b000000100000000011010101,
       24'b010010100010110011011111,
       24'b111110101111101011111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010101000011100111100010,
       24'b000000000000000011010110,
       24'b010111100100010111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b111001101110001011110101,
       24'b111101101111010111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111111111111101,
       24'b001111100001110011011110,
       24'b000000000000000011011001,
       24'b010011000011000011100001,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100010110111101011101011,
       24'b000000000000000011011000,
       24'b000101110000000011011100,
       24'b110101111101001011110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111011111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101001111001111111000,
       24'b101111111011110111110011,
       24'b110010001100011111110011,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b100100101000001011101000,
       24'b000000000000000011010101,
       24'b000000000000000011011011,
       24'b000101110000000011011001,
       24'b000010110000000011011010,
       24'b000000000000000011011001,
       24'b010010100010101011100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b010101000011101011100100,
       24'b000101010000100011011010,
       24'b001100010000111111011111,
       24'b000000000000000011011001,
       24'b101111011011001111110000,
       24'b111111111111111111111111,
       24'b101100111010011111101110,
       24'b000011010000000011011010,
       24'b001000110000000111011111,
       24'b000001010000000011011010,
       24'b010111100100001111100010,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010011000010111011100010,
       24'b000000000000000011010111,
       24'b011001100100110111100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010111100100000111011111,
       24'b000000000000000011010100,
       24'b011101000101111011101001,
       24'b111111111111111111111111,
       24'b100001010111001011101001,
       24'b000000000000000011010111,
       24'b001101100001001011011111,
       24'b111111001111110011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010011100000111110001,
       24'b000010010000000011011001,
       24'b000001100000000011011000,
       24'b110100011100110011110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101010001001101111110010,
       24'b000000000000000011010110,
       24'b001011100001000111011001,
       24'b111000011101110111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100010000111011011101001,
       24'b000000000000000011011000,
       24'b001100110001001111011111,
       24'b101011001001111111101110,
       24'b100010100111011111101010,
       24'b010010110011011011011111,
       24'b000010000000000011010101,
       24'b101110011010111111110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011011100101011111100100,
       24'b000000000000000011011000,
       24'b001010000000001111011110,
       24'b111100001110111011111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101101011010100111101111,
       24'b000001110000000011011000,
       24'b000010000000000011010111,
       24'b101000111001010111101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111011111110,
       24'b111111111111111111111010,
       24'b100000100111001111100111,
       24'b001010010001100011011011,
       24'b000000000000000011011000,
       24'b000000000000000011011001,
       24'b010010000011100111011110,
       24'b111001111110010111111000,
       24'b111111111111111111111111,
       24'b111101111111011011111010,
       24'b001010100000100111011100,
       24'b000010110000001011011010,
       24'b011000110100110011100110,
       24'b110101011100111111110010,
       24'b100011110111111111100111,
       24'b000010000000000011011100,
       24'b000000100000000011011000,
       24'b110010111100010111110001,
       24'b111111111111111111111111,
       24'b100001010111001011101001,
       24'b000000000000000011011000,
       24'b001010010000011011011111,
       24'b000000000000000011011010,
       24'b011000100100001111100100,
       24'b111111111111111111111111,
       24'b110000011011100011110100,
       24'b000010110000000011011100,
       24'b010000110010010111011111,
       24'b000111010000000011011011,
       24'b010000010010000111011110,
       24'b111110011111100111111010,
       24'b111111111111111111111111,
       24'b100000010110111011101000,
       24'b000000000000000011010110,
       24'b010001010010011111100001,
       24'b111111011111111011111100,
       24'b110011001100011011110010,
       24'b001010010001000011011110,
       24'b000000000000000011010110,
       24'b100000010110111111101001,
       24'b111111111111111111111111,
       24'b101100011010010011110000,
       24'b000001010000000011011001,
       24'b000101100000000011011010,
       24'b110011111100100111110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101101111011111111010,
       24'b001100010000101111011110,
       24'b000000000000000011010110,
       24'b100010110111101111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110110001101001111110100,
       24'b000010100000000011011010,
       24'b000001010000000011010111,
       24'b101111111011011011101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110111011001011110010,
       24'b000001100000000011011011,
       24'b000100110000000011011101,
       24'b000000000000000011010111,
       24'b000000000000000011010100,
       24'b000000000000000011010101,
       24'b000000000000000011010011,
       24'b100011010111101011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001101001100111101110,
       24'b000000000000000011011000,
       24'b000011100000000011011011,
       24'b110011011100011011110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011101110110011110110,
       24'b001011000000101111011010,
       24'b000000100000000111010111,
       24'b011110000110001011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100000010110111111100111,
       24'b000000000000000011010101,
       24'b000011110000000011011001,
       24'b001101110001001111011001,
       24'b000101000000000011011011,
       24'b000000000000000011011001,
       24'b010101010011010111100001,
       24'b111111111111111111111111,
       24'b111101101111011011111011,
       24'b001010000000010111100000,
       24'b000010100000010111010100,
       24'b101100101010100011101100,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b001011000000111011011111,
       24'b000001000000000111010111,
       24'b100111111001001011101010,
       24'b111111111111111111111111,
       24'b110000001011011111110000,
       24'b000010000000000011011001,
       24'b001100000000111111011100,
       24'b001000000000000011011100,
       24'b000110000000000011011100,
       24'b111111111111111111111011,
       24'b111001011110000111111000,
       24'b000001110000000011011011,
       24'b010110100100000011100000,
       24'b001101100001001111011111,
       24'b000010000000000011011011,
       24'b110100111100110111110100,
       24'b111111111111111111111111,
       24'b101010011001101111101111,
       24'b000000000000000011011000,
       24'b001011010000101111011110,
       24'b010000110010010111100000,
       24'b000011000000000011011010,
       24'b000000000000000011011001,
       24'b000100000000000011011001,
       24'b110111001101100011110100,
       24'b111111111111111111111111,
       24'b111000111101111111111000,
       24'b001010100000110011011100,
       24'b000010000000010011010111,
       24'b100100000111111111101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010010110010111011100010,
       24'b000011010000010011010110,
       24'b011100000101110111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111111111110,
       24'b111111111111111111111111,
       24'b111111101111111111111100,
       24'b001111010001100111011111,
       24'b000000000000000011010110,
       24'b011110110110100111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010001110010011110110,
       24'b000011010000000011010100,
       24'b000100000000000011011000,
       24'b010010010010110111100000,
       24'b011011010101101111100011,
       24'b100110111000111111100111,
       24'b110000111011111111101111,
       24'b111001101110001011111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110101001101000011110101,
       24'b000100110000000011011010,
       24'b000000000000000011011000,
       24'b100111011000111011101101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010001000010010011100010,
       24'b000000000000000011011001,
       24'b010110100011111011100010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110001111011111111011,
       24'b001011010000110011011110,
       24'b000000000000000011011011,
       24'b011010100101001011100100,
       24'b111010101110010111111001,
       24'b101001101001100011101101,
       24'b000001000000000011011011,
       24'b000010100000000011011010,
       24'b111001111110010111110110,
       24'b111111111111111111111111,
       24'b001110100001100111100001,
       24'b000000000000000011010110,
       24'b100000010110111111100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010101100011101011100001,
       24'b000000000000000011010111,
       24'b011001110100111111100101,
       24'b111111111111111111111111,
       24'b111010101110100011111000,
       24'b000101110000000011011011,
       24'b001111110001101011011101,
       24'b010100110011010011011111,
       24'b000000000000000011010111,
       24'b101111011011001011110000,
       24'b111111111111111111111010,
       24'b000001100000000011011001,
       24'b011000100100100111100010,
       24'b010111000100011011011110,
       24'b000000000000000011011000,
       24'b101001011001011011110000,
       24'b111111111111111111111111,
       24'b110011011100011011110011,
       24'b000100000000000011011001,
       24'b000111010000000011100000,
       24'b000001010000000011011011,
       24'b000011100000000011011010,
       24'b001110110010111011011101,
       24'b110010011011101111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b001110110001101011100000,
       24'b000000000000000011010101,
       24'b100011000111101011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101100110001011100111,
       24'b000001000000001011010111,
       24'b010000100010011011100000,
       24'b111111111111111111111011,
       24'b111110001111100011111001,
       24'b110011111100110111110011,
       24'b100110111001010111101010,
       24'b110101101101000011110011,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010110110100001011100011,
       24'b000000000000000011001111,
       24'b001010110000101011011100,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110101111101011111011,
       24'b101110111011000011101101,
       24'b110110011101101011110101,
       24'b111111111111111111111010,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101001111001111111011,
       24'b001011100000101011011110,
       24'b000000000000000011011000,
       24'b011010100101001111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010000101000011100110,
       24'b000000000000000011011001,
       24'b001100000001010111011100,
       24'b111011101110110111111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011111110111011110111,
       24'b001001100000001011011010,
       24'b000000000000000011011001,
       24'b101010111001111011101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b001010110000101011011101,
       24'b000000000000000011010001,
       24'b100010010111011111101010,
       24'b111111111111111111111111,
       24'b010111100100001111100011,
       24'b000000000000000011010110,
       24'b011000110100101011100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100000000110111111100110,
       24'b000000000000000011010111,
       24'b001110010001011011011111,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b001100110001000111011101,
       24'b000111100000011111011111,
       24'b100101011000100011101001,
       24'b000100100000000011011011,
       24'b010110000011100111100101,
       24'b111101011111011011110111,
       24'b000011110000000011011100,
       24'b011011100101011111101000,
       24'b100011000111110011100100,
       24'b000000010000000011010011,
       24'b011100110101111011100101,
       24'b111111111111111111111111,
       24'b111110101111101011111100,
       24'b001101100001000111011111,
       24'b000001010000000011011010,
       24'b010111010100101111100010,
       24'b110110001101011111110011,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010010101001011100010,
       24'b000110000000100111010110,
       24'b011010110101010111100001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011101010000111101111,
       24'b000001100000000011011001,
       24'b001001000000000111011111,
       24'b010110000011110111100001,
       24'b001101000001001011011110,
       24'b000010110000000011011011,
       24'b000000000000000011010000,
       24'b011101010110001011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101001101001100111101100,
       24'b010111100101101011100000,
       24'b101000111001010111101011,
       24'b111111111111111011111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011001100100111111100100,
       24'b000000000000000011011001,
       24'b010000010010001011100001,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100101101000011111101100,
       24'b000100100000010111011001,
       24'b001001000000100111011001,
       24'b101101101010101111110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111011111101,
       24'b010001110010101011100001,
       24'b000000000000000011010111,
       24'b011100000101101011100110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100100101110011100001,
       24'b010010100100001111011011,
       24'b101110101011000011110001,
       24'b111111111111111111111111,
       24'b100011010111110011101011,
       24'b000000000000000011010111,
       24'b001100110001000011011100,
       24'b111100001111000011111000,
       24'b111111111111111111111111,
       24'b101101101010110111110000,
       24'b000000000000000011011000,
       24'b000110010000000011011101,
       24'b111001011110001111111001,
       24'b111111111111111111111111,
       24'b011011000101010111100110,
       24'b000000000000000011010101,
       24'b101001011001011111101010,
       24'b011010100100111011100101,
       24'b000000000000000011011000,
       24'b101111111011011011110000,
       24'b010000010010000011100001,
       24'b011101000110000011101000,
       24'b101001101001011111101111,
       24'b000001000000000011010101,
       24'b010100010011010111011100,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b011000010100100011100101,
       24'b000000000000000011010101,
       24'b011010100101000111100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100111011001000011101011,
       24'b000101110000101111011001,
       24'b001001000000000011011110,
       24'b110110111101010111110010,
       24'b110001001011110011110000,
       24'b100001000111101011101000,
       24'b010101110100111111100001,
       24'b111010111110100111111000,
       24'b111100001110111011111010,
       24'b000100000000000011011011,
       24'b000000000000000011011010,
       24'b000000000000000011010101,
       24'b000000000000000011011000,
       24'b000101100000000011011100,
       24'b001001100010001011011011,
       24'b100111011000111111101001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111111111111100,
       24'b110110011101011011110101,
       24'b101001111001111011101011,
       24'b011111010110111011101000,
       24'b001110100010010111100001,
       24'b001001010000110111011011,
       24'b001011100000111011011011,
       24'b110101011101000011110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110010111100001111110011,
       24'b001001000000001011011001,
       24'b000111000001000011010111,
       24'b100101111000011011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011100000101100111100111,
       24'b000000000000000011010111,
       24'b010001100010011011100010,
       24'b111111111111111111111110,
       24'b111111111111111111111110,
       24'b111111111111110111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110000111011101011110010,
       24'b000010010000000011011001,
       24'b000001100000000011011010,
       24'b110000101011100111110010,
       24'b111111111111111111111111,
       24'b110101111101001111110111,
       24'b000100000000000011011100,
       24'b000001100000000011011001,
       24'b101111101011010011110001,
       24'b111111111111111111111111,
       24'b100100011000000011101101,
       24'b000010000000001011010100,
       24'b101110101011000011101011,
       24'b101101001010100111101111,
       24'b000000000000000011010111,
       24'b011100100101101011100100,
       24'b010011000010111011011110,
       24'b011010100101010011100111,
       24'b110000101011100111110000,
       24'b000000000000000011011010,
       24'b000111100000000011011101,
       24'b111010101110011011111000,
       24'b111111111111111111111111,
       24'b100000000110111011101001,
       24'b000000000000000011010111,
       24'b001110110001011111100000,
       24'b111111011111110011111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001011011111011110010,
       24'b000001000000000011011001,
       24'b001000000000000011011110,
       24'b001001010000000111011100,
       24'b000000000000000011011000,
       24'b000000000000000011010110,
       24'b000000000000000011001111,
       24'b101000011001010011101101,
       24'b111111111111111111111110,
       24'b001111000001110111011011,
       24'b010001100011101111011111,
       24'b100010100111110111101000,
       24'b101111011011011011110001,
       24'b110111001101110011110101,
       24'b111111111111111111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111100,
       24'b111001101110011011111000,
       24'b101110101011010011110000,
       24'b100000110111011111100111,
       24'b010101110100001011100001,
       24'b001110010001111111011111,
       24'b000111000000000011011100,
       24'b000000000000000011011001,
       24'b000000000000000011011000,
       24'b000000000000000011011011,
       24'b000001010000000011011011,
       24'b001000100000010011010101,
       24'b110001011011110011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111110011111100,
       24'b001100100001000111011111,
       24'b000000000000000011010111,
       24'b011100100101110011100111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100100111000001111101010,
       24'b000000000000000011011000,
       24'b001010010000010111011101,
       24'b111011111110111111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111100111111000111111001,
       24'b001010110000100011011101,
       24'b000000000000000011010111,
       24'b101000011001001111101111,
       24'b111111111111111111111111,
       24'b111110001111100011111011,
       24'b001100100000110011011111,
       24'b000000000000000011010110,
       24'b100001110111010111101001,
       24'b111111111111111111111111,
       24'b101101101010110011110000,
       24'b000000010000000011011000,
       24'b011000000100000011100101,
       24'b111000101101111111110101,
       24'b000111110000001011011111,
       24'b000111100000000011011100,
       24'b000111010000011011011010,
       24'b011000010100011111101000,
       24'b111000111110001011110101,
       24'b001001000000011011011101,
       24'b000011110000000011011001,
       24'b110001101011110111110010,
       24'b111111111111111111111111,
       24'b101011001001111111101110,
       24'b000000000000000011011010,
       24'b000100110000000011011011,
       24'b110110101101010011110110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010011110011011110110,
       24'b000001010000000011011000,
       24'b000000000000000011010101,
       24'b000001010000000011011000,
       24'b001010010000100111011101,
       24'b010011000011010011100001,
       24'b011010010110001111100010,
       24'b110010001100001011110011,
       24'b111111111111111111111111,
       24'b111101101111010111111000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b111001101110011111110111,
       24'b110010001100001111110010,
       24'b100110101001000011101010,
       24'b011010000101010111100100,
       24'b010001010010110111100001,
       24'b001010110000110011011110,
       24'b000010000000000011011001,
       24'b000000000000000011011000,
       24'b000000000000000011011001,
       24'b000000000000000011011001,
       24'b000000000000000011010111,
       24'b000000110000000011010110,
       24'b000111000000000011011011,
       24'b001110110001111111011111,
       24'b010011000100001011100000,
       24'b101011011010000111101010,
       24'b111111111111111111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b010100110011100011100011,
       24'b000000000000000011011001,
       24'b010001000010010111011101,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110001101011111111110010,
       24'b000010100000000011011001,
       24'b000001000000000011011001,
       24'b101110111011001111110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010010010010101011100010,
       24'b000000000000000011010111,
       24'b011101110110001011101000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011000010100011111100100,
       24'b000000000000000011010111,
       24'b010100110011011111100010,
       24'b111111111111111111111111,
       24'b111100001110111111111001,
       24'b000110010000000111011011,
       24'b000010000000000011011101,
       24'b111111001111110111111000,
       24'b100001010110111111101010,
       24'b000000000000000011011001,
       24'b000010110000000011011011,
       24'b010010010010110011100101,
       24'b111111111111111111111011,
       24'b010101110011100011100011,
       24'b000000100000000011010101,
       24'b100100101000001011101010,
       24'b111111111111111111111111,
       24'b111000001101110011110111,
       24'b001001000000101111011100,
       24'b000001110000000011010101,
       24'b100111111001000111101011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111001111110111111010,
       24'b100000100110110011100101,
       24'b100001111000000111100111,
       24'b110000111011111111110010,
       24'b111011111111000011111010,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111011111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111011111110111011110101,
       24'b110000111011110011110000,
       24'b101000011001011111101101,
       24'b011110100110100111100110,
       24'b010010000011000111011110,
       24'b001001010000100011011010,
       24'b000100000000000011011010,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000110010000000011011010,
       24'b001110110010000011011100,
       24'b010110100100011011100010,
       24'b011111010110111111100110,
       24'b101010101010000111101100,
       24'b110110011101100011110101,
       24'b111111001111111011111010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011111110110111011101000,
       24'b000000000000000011011000,
       24'b001000010000001011011010,
       24'b111001001110000111110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111101011111010111111010,
       24'b001011100000110011011110,
       24'b000000000000000011011000,
       24'b100011000111100111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111011111011,
       24'b111110011111100111111011,
       24'b111111111111111111111111,
       24'b011100000101101111100101,
       24'b000000010000000011010111,
       24'b010001000010010111011111,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b100100101000000111101011,
       24'b000000010000000011011001,
       24'b001010110000100011011101,
       24'b111101101111010011111011,
       24'b111111111111111111111111,
       24'b010011100010110011100011,
       24'b000000000000000011010110,
       24'b110111111101101111110111,
       24'b111010001110010111110111,
       24'b000000000000000011010111,
       24'b000011110000000011011111,
       24'b010000110010011111100000,
       24'b111111111111111111111101,
       24'b011110010110010011101010,
       24'b000000000000000011010110,
       24'b010110010100000011100100,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b001011000000100111011010,
       24'b000000000000000011001110,
       24'b011010110101010011100100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111010,
       24'b111001101110001011110010,
       24'b110000111011110011101001,
       24'b100000100111010011101000,
       24'b010100010100000111100011,
       24'b001111110010001111011001,
       24'b000110010000000011011000,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b000100110000000011011010,
       24'b001010010000110011011011,
       24'b010100000011110011100000,
       24'b011111110111000011100111,
       24'b101001011001110011101100,
       24'b110001111100001111110010,
       24'b111101001111010111111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110001010110111110000,
       24'b000000010000000011011001,
       24'b000000110000000011011010,
       24'b101111101011010011110001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010101000011101111100001,
       24'b000000010000000011010110,
       24'b011010110101010011100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100100001000000111101000,
       24'b001000010001111011010111,
       24'b011101110110001011100101,
       24'b111111111111111111111111,
       24'b101011001010000111101100,
       24'b000000110000000011010110,
       24'b000111110000000011011101,
       24'b111011011110101111111001,
       24'b111111111111111111111111,
       24'b101111111011011011110010,
       24'b000001100000000011011001,
       24'b000100100000000011011100,
       24'b110011111100100111110100,
       24'b111111111111111111111111,
       24'b011100110101110111100111,
       24'b000000000000000011010010,
       24'b100011000111110011101011,
       24'b111111111111111111111111,
       24'b001111000001101111011111,
       24'b000000000000000011011100,
       24'b001010110000101011011101,
       24'b111111111111111111111111,
       24'b100110111000111011101011,
       24'b000000000000000011001110,
       24'b001010110000101011011100,
       24'b111111001111110111111100,
       24'b111111111111111111111111,
       24'b101000111001011011101010,
       24'b101000011010000111101011,
       24'b110111101101100111110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111001101110010011110100,
       24'b101100011010101011101101,
       24'b100000110111001111100111,
       24'b010010110011001011100011,
       24'b010000010010011011011111,
       24'b001111010010000011010110,
       24'b001001100000010011010011,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b001001000000000111011100,
       24'b001001110000100011010111,
       24'b000000100000000011011000,
       24'b000111010000000011011100,
       24'b001111100010011011011111,
       24'b011011010101110111100100,
       24'b101000111001011111101011,
       24'b110010111100100111110010,
       24'b111010101110110011111000,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110111011101100011110111,
       24'b000111110000000111011011,
       24'b000000000000000011010111,
       24'b100010010111011111101010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101010101111111100110,
       24'b000000000000000011011000,
       24'b010000110010000111100000,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b011110110110011011101000,
       24'b000000000000000011010011,
       24'b001110110001101011011111,
       24'b111111111111111111111111,
       24'b111000001101110111110110,
       24'b000001100000000011011001,
       24'b000000110000000011011010,
       24'b110000011011100111110000,
       24'b111111111111111111111111,
       24'b110010111100010011110001,
       24'b000001100000000011010111,
       24'b000010000000000011011011,
       24'b110001001011110011110100,
       24'b111111111111111111111111,
       24'b101011001010000111101010,
       24'b000000000000000011010100,
       24'b001101000001001111100001,
       24'b111111111111111111111111,
       24'b100011100111101111101010,
       24'b000000000000000011010001,
       24'b001011010000101111011010,
       24'b111101111111011111111100,
       24'b111000101101111011110101,
       24'b100011111000100111101000,
       24'b110010011100001011110011,
       24'b111111011111110011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b111000111110000111110110,
       24'b110000111011111011110011,
       24'b100101111000100111101011,
       24'b011000110101000111100010,
       24'b010000100010100111011111,
       24'b000111110000000011011100,
       24'b000010100000000011011000,
       24'b000110110000000011010101,
       24'b000011100000000011010110,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000010000000011011001,
       24'b001001010000000111011011,
       24'b010010100011000111011110,
       24'b011001010101010011100001,
       24'b100101111000101011101000,
       24'b101110111011011011110010,
       24'b110111011101110111110110,
       24'b111111111111111111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110101111101011111011,
       24'b001110110001101011011101,
       24'b000000000000000011011001,
       24'b010100100011011111100010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101011001010000111101100,
       24'b000000000000000011011000,
       24'b000110010000000011011011,
       24'b111001001110000111110111,
       24'b111111111111111111111111,
       24'b110101111101000011110110,
       24'b000001010000000011011010,
       24'b000110010000000011011011,
       24'b111100011111000111111001,
       24'b111111111111111111111110,
       24'b001100010000110011011101,
       24'b000000000000000011011010,
       24'b001111100001111011011111,
       24'b100100010111111111101000,
       24'b010011010010111011100010,
       24'b000000000000000011011100,
       24'b000110000000000011011010,
       24'b111010101110011011111001,
       24'b111111111111111111111111,
       24'b110011111100100011110011,
       24'b000000000000000011010100,
       24'b010011100011001111011110,
       24'b111111011111110111111100,
       24'b111011101110110011111001,
       24'b101100011010110111101100,
       24'b111010111110101011110101,
       24'b111110101111101011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111011101110111011111001,
       24'b110000101011111011110010,
       24'b100111101001010011101101,
       24'b011101010110010111100110,
       24'b010010110011011011011101,
       24'b001001010000100111011101,
       24'b000011000000000011011010,
       24'b000000000000000011010111,
       24'b000000000000000011011000,
       24'b000000000000000011011011,
       24'b000000000000000011011001,
       24'b000010100000000011010111,
       24'b001101010001111111010011,
       24'b100000100111000011010111,
       24'b011010010101011011100101,
       24'b011111000110110111101001,
       24'b101010001010000111101110,
       24'b111000011101111111110101,
       24'b111111111111111111111100,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011010100101001111100110,
       24'b000000000000000011011000,
       24'b001011010000100111011110,
       24'b111100111111001111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111001001110000111110110,
       24'b001000110000100111011001,
       24'b000000000000000011011001,
       24'b101010011001111011101101,
       24'b111111111111111111111111,
       24'b110010111100001111110010,
       24'b000101100000001011011100,
       24'b001001010000101011011011,
       24'b110101011100111111110101,
       24'b111111111111111111111111,
       24'b101101011010101111101111,
       24'b000000000000000011010110,
       24'b000000000000000011011001,
       24'b000000000000000011010111,
       24'b000000000000000011010101,
       24'b000001000000000011011000,
       24'b101011011010000011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111101011111010011111010,
       24'b110110111101001111110010,
       24'b111111011111111011111000,
       24'b111111101111111011111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111001111110011111010,
       24'b110101101101001011110010,
       24'b101000001001100011101010,
       24'b011110000110100111101000,
       24'b010101100011111111100010,
       24'b001011010001000111011100,
       24'b000011100000000011011000,
       24'b000000000000000011011000,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011011001,
       24'b000010100000000011011010,
       24'b001001100000100111011010,
       24'b010011110011101011011111,
       24'b100011010111111011100110,
       24'b101011011010001111101100,
       24'b110000011011110011110010,
       24'b111110101111110011111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110011000100111101100,
       24'b000000000000000011011000,
       24'b000100110000000011011100,
       24'b110100011100100111110100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b010001110010010111100000,
       24'b000000000000000011011011,
       24'b001101110001001111100000,
       24'b011101110110000111100100,
       24'b001110010001011011011111,
       24'b000000100000000011011010,
       24'b010010010010111011011110,
       24'b111011111110110011111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111011010110111101111,
       24'b010110100101000011100010,
       24'b010110000100010011011110,
       24'b011111110111100111100110,
       24'b110011111100010011110010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b111000001110000111110111,
       24'b101100111010110111101110,
       24'b100001010111100011100111,
       24'b010111010100110111100100,
       24'b010111000100010011011010,
       24'b001110010001101111010101,
       24'b000000000000000011011010,
       24'b000000000000000011011011,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000011000000000011011011,
       24'b001000010000000111011011,
       24'b010000000010011011011101,
       24'b011100000101111111100011,
       24'b100111101001001111101011,
       24'b101111111011100111110010,
       24'b111010011110101011110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101110011010111011110010,
       24'b000010000000000011011010,
       24'b000000010000000011011000,
       24'b101001111001101011101110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b101111101011010111110001,
       24'b000001000000000011010111,
       24'b000000000000000011010111,
       24'b000000000000000011010101,
       24'b000000000000000011010101,
       24'b000100000000010111011000,
       24'b101110011011000011110000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111010,
       24'b111000001110000111110101,
       24'b110001111100000111101111,
       24'b100100011000011011101000,
       24'b011010000101010111100011,
       24'b010001100010101111011111,
       24'b000111100000000111011011,
       24'b000001010000000011010110,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000011110000000011010101,
       24'b000000000000000011010110,
       24'b000001100000000011011000,
       24'b001000100000000111011011,
       24'b001111100010011011100000,
       24'b011000000100110011100011,
       24'b100100111000010111101000,
       24'b110000001011101011110000,
       24'b111000001110000011110101,
       24'b111111111111111111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111010011110010111111001,
       24'b001001010000000011011100,
       24'b000000000000000011011000,
       24'b011011110101101011100101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110011101100000111110001,
       24'b011010100110010011100100,
       24'b011010000101101111100101,
       24'b100001111000000011100111,
       24'b111010011110000011110101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111101,
       24'b111011001110110011110101,
       24'b101110111011010111101111,
       24'b100110101001000011101100,
       24'b011101100110010011100110,
       24'b010001010010110011011110,
       24'b001000010000001111011011,
       24'b000111000000000011011000,
       24'b000010110000000011010111,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b000000000000000011011000,
       24'b000110110000000011011001,
       24'b010000000010011011011101,
       24'b010110110100100011100100,
       24'b100000010111001011101001,
       24'b101100101010110111101011,
       24'b111000001101111111110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b010011010010111111100010,
       24'b000000000000000011011001,
       24'b010010010010101011100010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111110011111101011111011,
       24'b110011011100101011110000,
       24'b101010001010000011101100,
       24'b100001000111010111100111,
       24'b010100110011110011100000,
       24'b001001100000101011011011,
       24'b000110010000000011011000,
       24'b000000010000000011010111,
       24'b000000000000000011011011,
       24'b000101000000000011011100,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000100100000000011011001,
       24'b001100000001010011011010,
       24'b010101110100000111100010,
       24'b011101110110100011100111,
       24'b101000001001010111101100,
       24'b110100001100111011110010,
       24'b111110111111110111111001,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b011101000101111111100111,
       24'b000000000000000011011000,
       24'b001010100000011011011110,
       24'b111100001110111111111000,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111101111111111111100,
       24'b110111111101110111110110,
       24'b101011101010010111101101,
       24'b011111110111000111101000,
       24'b011000110100111011100100,
       24'b001110100001111011011101,
       24'b000110110000000011010111,
       24'b000001000000000011011001,
       24'b000000000000000011011001,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000001110000000011010110,
       24'b000100010000000011011000,
       24'b001000010000001111011100,
       24'b010011000011011111011111,
       24'b011101010110010011100101,
       24'b100111001001001011101101,
       24'b101111101011100111110001,
       24'b111011001110110011110111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110011000101011101100,
       24'b000000000000000011011000,
       24'b000010000000000011011001,
       24'b101110111011001111101111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b110111111101111011110111,
       24'b110001001011110111110010,
       24'b100011111000001111101001,
       24'b011000000100110111100010,
       24'b001111000010001011011110,
       24'b000111110000000011011011,
       24'b000010000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011011,
       24'b000001100000000011011001,
       24'b001000010000001111011011,
       24'b010100110011100111011101,
       24'b011010100101100011100001,
       24'b100100111000011011101011,
       24'b110000011011110011110100,
       24'b111000011110000111110111,
       24'b111111111111111111111011,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b110100101100110011110011,
       24'b000000000000000011010101,
       24'b000000000000000011010111,
       24'b100101001000001111101100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111100,
       24'b111011001110110111110111,
       24'b110010111100100011110011,
       24'b101000011001010111101011,
       24'b011011010101111011100100,
       24'b001111100010011111011110,
       24'b001000000000001011011100,
       24'b000100100000000011011000,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000000000000000011011010,
       24'b000000000000000011011001,
       24'b000001010000000011010111,
       24'b001000000000000011011010,
       24'b001101100001101111011111,
       24'b010100110011110111100001,
       24'b100000000111000111100110,
       24'b101100111010110111101110,
       24'b111000101110001011110101,
       24'b111111111111111111111010,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b101101111010100111101110,
       24'b000000000000000011010110,
       24'b010110110100011111100100,
       24'b110110001101000011110100,
       24'b101010001010000011101111,
       24'b100000100111001111101000,
       24'b010100010011100111100000,
       24'b001000110000010011011011,
       24'b000101000000000011011010,
       24'b000001010000000011011001,
       24'b000000000000000011011011,
       24'b000000000000000011011010,
       24'b000000000000000011011000,
       24'b000000000000000011011001,
       24'b000011010000000011011011,
       24'b001011110001000011011011,
       24'b010110010100001111100010,
       24'b011111000110101011100110,
       24'b101000011001011111101010,
       24'b110100111101000011110100,
       24'b111110101111110011111010,
       24'b111111111111111111111110,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111110,
       24'b100111101000100111101011,
       24'b000000000000000011010110,
       24'b000011100000000011011010,
       24'b000000110000000011011011,
       24'b000000000000000011011000,
       24'b000000000000000011011010,
       24'b000100000000000011011100,
       24'b000000000000000011011000,
       24'b000101110000000011011011,
       24'b001000100000011011011010,
       24'b010010100011001111011101,
       24'b011111000110110011100110,
       24'b100111101001010111101100,
       24'b110000101011110111110000,
       24'b111100001111000011110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111011111110011111110,
       24'b011110010110010011100101,
       24'b100111111001001111101011,
       24'b110011111100101011110010,
       24'b000010010000000011011000,
       24'b000000000000000011010110,
       24'b001001010000011111011011,
       24'b010010110011011011100000,
       24'b011110100110111011100100,
       24'b100110001000110111101010,
       24'b110000011011110111110001,
       24'b111001011110011011110110,
       24'b111111111111111111111101,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b100110011000100111101101,
       24'b000100110000011011010101,
       24'b111101111111010111110111,
       24'b110001011011101111110001,
       24'b101001111010001111101100,
       24'b111001011110010111110111,
       24'b111111111111111111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111011,
       24'b111100001111001011110111,
       24'b111100111111000111111100,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
       24'b111111111111111111111111,
};

// define maze param
// see maze.txt
localparam [0:4][4:0] maze = {5'b00000, 5'b10101, 5'b10100, 5'b10011, 5'b00111};
localparam [0:5][4:0] hor_wall = {5'b11111, 5'b10101, 5'b00001, 5'b00111, 5'b10100, 5'b11111};
localparam [0:5][4:0] ver_wall = {5'b11111, 5'b00010, 5'b01110, 5'b10110, 5'b01110, 5'b11111};
//reg [2:0] pos[1:0] = {1'b0, 1'b0};

//define camera param
localparam width = 10'd800;
localparam height = 10'd600;
localparam unit_size = 8'd64;
reg [1:0] dir;
localparam U = 2'd0;
localparam L = 2'd1;
localparam D = 2'd2;
localparam R = 2'd3;
reg [2:0] x;
reg [2:0] y;

// define state
reg [3:0] state = 4'b0000;
localparam STILL = 4'b0001;
localparam INIT_CAM = 4'b0010;
localparam DRAW = 4'b0011;

reg [3:0] enter_state = 4'b0100;
localparam NONE = 4'b0000;
localparam COVER_PHASE1 = 4'b0100;
localparam COVER_PHASE2 = 4'b0101;
localparam FINAL_PHASE = 4'b0110;
localparam ENTER_PHASE1 = 4'b0001;
localparam ENTER_PHASE2 = 4'b0010;
localparam ENTER_PHASE3 = 4'b0011;

reg[7:0] grad_cnt = 8'd0;
reg[16:0] grad_rate = 17'd0;

// define movement signal
reg [3:0] draw_mode = 4'b0000; // 01 move 10 left 11 right
localparam MOVE = 4'b0001;
localparam LEFT = 4'b0010;
localparam RIGHT = 4'b0011;
localparam DARKEN = 4'b0100;
localparam UP = 4'b0101;
localparam DOWN = 4'b0110;

reg [8:0] pip_en; // 使能 拉低有效
reg [9:0] px[8:0]; // 像素点x
reg [9:0] py[8:0]; // 像素点y

// LED
// assign leds[1:0] = move_data;
// assign leds[2] = wr_en;
// assign leds[15:3] = 12'd0;
// assign leds[31:16] = ~(dip_sw);

wire signal;
wire move_data_addtion;

ps2_controller u_ps2_controller(
    .clk(clk_ps2), // 50MHz
    .rst(reset_btn),
    .ps2_clk(ps2_clock),
    .ps2_data(ps2_data),
    .data(move_data),
    .signal(signal),
    .move_data_addtion(move_data_addtion)
);

wire [3:0] move_data;
reg move_en = 0;

reg [31:0] offset_reg = 1'b0;
wire rd_addr_offset;
wire wr_addr_offset;

assign rd_addr_offset = offset_reg[0];
assign wr_addr_offset = ~offset_reg[0];

reg wr_en = 1'b0;
reg [18:0] wr_addr = 19'b0;
wire [31:0] wr_data;
reg [7:0] image_cnt = 8'd0;
reg signed [9:0] center_x = unit_size >> 1;
reg signed [9:0] center_y = unit_size >> 1;
reg signed [9:0] center_z = 120;
reg [8:0] center_angle = 9'd180;
localparam signed [0:359][9:0] Dir_x = {
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000010,
    10'b1000000011,
    10'b1000000100,
    10'b1000000101,
    10'b1000000110,
    10'b1000001000,
    10'b1000001001,
    10'b1000001011,
    10'b1000001101,
    10'b1000001111,
    10'b1000010001,
    10'b1000010100,
    10'b1000010110,
    10'b1000011001,
    10'b1000011100,
    10'b1000011111,
    10'b1000100010,
    10'b1000100101,
    10'b1000101001,
    10'b1000101100,
    10'b1000110000,
    10'b1000110100,
    10'b1000111000,
    10'b1000111100,
    10'b1001000000,
    10'b1001000101,
    10'b1001001001,
    10'b1001001110,
    10'b1001010011,
    10'b1001011000,
    10'b1001011101,
    10'b1001100010,
    10'b1001100111,
    10'b1001101101,
    10'b1001110010,
    10'b1001111000,
    10'b1001111110,
    10'b1010000100,
    10'b1010001010,
    10'b1010010000,
    10'b1010010110,
    10'b1010011100,
    10'b1010100011,
    10'b1010101001,
    10'b1010110000,
    10'b1010110111,
    10'b1010111110,
    10'b1011000101,
    10'b1011001100,
    10'b1011010011,
    10'b1011011010,
    10'b1011100010,
    10'b1011101001,
    10'b1011110001,
    10'b1011111000,
    10'b1100000000,
    10'b1100001000,
    10'b1100010000,
    10'b1100011000,
    10'b1100100000,
    10'b1100101000,
    10'b1100110000,
    10'b1100111000,
    10'b1101000000,
    10'b1101001001,
    10'b1101010001,
    10'b1101011001,
    10'b1101100010,
    10'b1101101010,
    10'b1101110011,
    10'b1101111011,
    10'b1110000100,
    10'b1110001101,
    10'b1110010110,
    10'b1110011110,
    10'b1110100111,
    10'b1110110000,
    10'b1110111001,
    10'b1111000010,
    10'b1111001010,
    10'b1111010011,
    10'b1111011100,
    10'b1111100101,
    10'b1111101110,
    10'b1111110111,
    10'b0000000000,
    10'b0000001001,
    10'b0000010010,
    10'b0000011011,
    10'b0000100100,
    10'b0000101101,
    10'b0000110110,
    10'b0000111110,
    10'b0001000111,
    10'b0001010000,
    10'b0001011001,
    10'b0001100010,
    10'b0001101010,
    10'b0001110011,
    10'b0001111100,
    10'b0010000101,
    10'b0010001101,
    10'b0010010110,
    10'b0010011110,
    10'b0010100111,
    10'b0010101111,
    10'b0010110111,
    10'b0011000000,
    10'b0011001000,
    10'b0011010000,
    10'b0011011000,
    10'b0011100000,
    10'b0011101000,
    10'b0011110000,
    10'b0011111000,
    10'b0100000000,
    10'b0100001000,
    10'b0100001111,
    10'b0100010111,
    10'b0100011110,
    10'b0100100110,
    10'b0100101101,
    10'b0100110100,
    10'b0100111011,
    10'b0101000010,
    10'b0101001001,
    10'b0101010000,
    10'b0101010111,
    10'b0101011101,
    10'b0101100100,
    10'b0101101010,
    10'b0101110000,
    10'b0101110110,
    10'b0101111100,
    10'b0110000010,
    10'b0110001000,
    10'b0110001110,
    10'b0110010011,
    10'b0110011001,
    10'b0110011110,
    10'b0110100011,
    10'b0110101000,
    10'b0110101101,
    10'b0110110010,
    10'b0110110111,
    10'b0110111011,
    10'b0111000000,
    10'b0111000100,
    10'b0111001000,
    10'b0111001100,
    10'b0111010000,
    10'b0111010100,
    10'b0111010111,
    10'b0111011011,
    10'b0111011110,
    10'b0111100001,
    10'b0111100100,
    10'b0111100111,
    10'b0111101010,
    10'b0111101100,
    10'b0111101111,
    10'b0111110001,
    10'b0111110011,
    10'b0111110101,
    10'b0111110111,
    10'b0111111000,
    10'b0111111010,
    10'b0111111011,
    10'b0111111100,
    10'b0111111101,
    10'b0111111110,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111110,
    10'b0111111101,
    10'b0111111100,
    10'b0111111011,
    10'b0111111010,
    10'b0111111000,
    10'b0111110111,
    10'b0111110101,
    10'b0111110011,
    10'b0111110001,
    10'b0111101111,
    10'b0111101100,
    10'b0111101010,
    10'b0111100111,
    10'b0111100100,
    10'b0111100001,
    10'b0111011110,
    10'b0111011011,
    10'b0111010111,
    10'b0111010100,
    10'b0111010000,
    10'b0111001100,
    10'b0111001000,
    10'b0111000100,
    10'b0111000000,
    10'b0110111011,
    10'b0110110111,
    10'b0110110010,
    10'b0110101101,
    10'b0110101000,
    10'b0110100011,
    10'b0110011110,
    10'b0110011001,
    10'b0110010011,
    10'b0110001110,
    10'b0110001000,
    10'b0110000010,
    10'b0101111100,
    10'b0101110110,
    10'b0101110000,
    10'b0101101010,
    10'b0101100100,
    10'b0101011101,
    10'b0101010111,
    10'b0101010000,
    10'b0101001001,
    10'b0101000010,
    10'b0100111011,
    10'b0100110100,
    10'b0100101101,
    10'b0100100110,
    10'b0100011110,
    10'b0100010111,
    10'b0100001111,
    10'b0100001000,
    10'b0100000000,
    10'b0011111000,
    10'b0011110000,
    10'b0011101000,
    10'b0011100000,
    10'b0011011000,
    10'b0011010000,
    10'b0011001000,
    10'b0011000000,
    10'b0010110111,
    10'b0010101111,
    10'b0010100111,
    10'b0010011110,
    10'b0010010110,
    10'b0010001101,
    10'b0010000101,
    10'b0001111100,
    10'b0001110011,
    10'b0001101010,
    10'b0001100010,
    10'b0001011001,
    10'b0001010000,
    10'b0001000111,
    10'b0000111110,
    10'b0000110110,
    10'b0000101101,
    10'b0000100100,
    10'b0000011011,
    10'b0000010010,
    10'b0000001001,
    10'b0000000000,
    10'b1111110111,
    10'b1111101110,
    10'b1111100101,
    10'b1111011100,
    10'b1111010011,
    10'b1111001010,
    10'b1111000010,
    10'b1110111001,
    10'b1110110000,
    10'b1110100111,
    10'b1110011110,
    10'b1110010110,
    10'b1110001101,
    10'b1110000100,
    10'b1101111011,
    10'b1101110011,
    10'b1101101010,
    10'b1101100010,
    10'b1101011001,
    10'b1101010001,
    10'b1101001001,
    10'b1101000000,
    10'b1100111000,
    10'b1100110000,
    10'b1100101000,
    10'b1100100000,
    10'b1100011000,
    10'b1100010000,
    10'b1100001000,
    10'b1100000000,
    10'b1011111000,
    10'b1011110001,
    10'b1011101001,
    10'b1011100010,
    10'b1011011010,
    10'b1011010011,
    10'b1011001100,
    10'b1011000101,
    10'b1010111110,
    10'b1010110111,
    10'b1010110000,
    10'b1010101001,
    10'b1010100011,
    10'b1010011100,
    10'b1010010110,
    10'b1010010000,
    10'b1010001010,
    10'b1010000100,
    10'b1001111110,
    10'b1001111000,
    10'b1001110010,
    10'b1001101101,
    10'b1001100111,
    10'b1001100010,
    10'b1001011101,
    10'b1001011000,
    10'b1001010011,
    10'b1001001110,
    10'b1001001001,
    10'b1001000101,
    10'b1001000000,
    10'b1000111100,
    10'b1000111000,
    10'b1000110100,
    10'b1000110000,
    10'b1000101100,
    10'b1000101001,
    10'b1000100101,
    10'b1000100010,
    10'b1000011111,
    10'b1000011100,
    10'b1000011001,
    10'b1000010110,
    10'b1000010100,
    10'b1000010001,
    10'b1000001111,
    10'b1000001101,
    10'b1000001011,
    10'b1000001001,
    10'b1000001000,
    10'b1000000110,
    10'b1000000101,
    10'b1000000100,
    10'b1000000011,
    10'b1000000010,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001
};
localparam signed [0:359][9:0] Dir_y = {
    10'b0000000000,
    10'b0000001001,
    10'b0000010010,
    10'b0000011011,
    10'b0000100100,
    10'b0000101101,
    10'b0000110110,
    10'b0000111110,
    10'b0001000111,
    10'b0001010000,
    10'b0001011001,
    10'b0001100010,
    10'b0001101010,
    10'b0001110011,
    10'b0001111100,
    10'b0010000101,
    10'b0010001101,
    10'b0010010110,
    10'b0010011110,
    10'b0010100111,
    10'b0010101111,
    10'b0010110111,
    10'b0011000000,
    10'b0011001000,
    10'b0011010000,
    10'b0011011000,
    10'b0011100000,
    10'b0011101000,
    10'b0011110000,
    10'b0011111000,
    10'b0100000000,
    10'b0100001000,
    10'b0100001111,
    10'b0100010111,
    10'b0100011110,
    10'b0100100110,
    10'b0100101101,
    10'b0100110100,
    10'b0100111011,
    10'b0101000010,
    10'b0101001001,
    10'b0101010000,
    10'b0101010111,
    10'b0101011101,
    10'b0101100100,
    10'b0101101010,
    10'b0101110000,
    10'b0101110110,
    10'b0101111100,
    10'b0110000010,
    10'b0110001000,
    10'b0110001110,
    10'b0110010011,
    10'b0110011001,
    10'b0110011110,
    10'b0110100011,
    10'b0110101000,
    10'b0110101101,
    10'b0110110010,
    10'b0110110111,
    10'b0110111011,
    10'b0111000000,
    10'b0111000100,
    10'b0111001000,
    10'b0111001100,
    10'b0111010000,
    10'b0111010100,
    10'b0111010111,
    10'b0111011011,
    10'b0111011110,
    10'b0111100001,
    10'b0111100100,
    10'b0111100111,
    10'b0111101010,
    10'b0111101100,
    10'b0111101111,
    10'b0111110001,
    10'b0111110011,
    10'b0111110101,
    10'b0111110111,
    10'b0111111000,
    10'b0111111010,
    10'b0111111011,
    10'b0111111100,
    10'b0111111101,
    10'b0111111110,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111111,
    10'b0111111110,
    10'b0111111101,
    10'b0111111100,
    10'b0111111011,
    10'b0111111010,
    10'b0111111000,
    10'b0111110111,
    10'b0111110101,
    10'b0111110011,
    10'b0111110001,
    10'b0111101111,
    10'b0111101100,
    10'b0111101010,
    10'b0111100111,
    10'b0111100100,
    10'b0111100001,
    10'b0111011110,
    10'b0111011011,
    10'b0111010111,
    10'b0111010100,
    10'b0111010000,
    10'b0111001100,
    10'b0111001000,
    10'b0111000100,
    10'b0111000000,
    10'b0110111011,
    10'b0110110111,
    10'b0110110010,
    10'b0110101101,
    10'b0110101000,
    10'b0110100011,
    10'b0110011110,
    10'b0110011001,
    10'b0110010011,
    10'b0110001110,
    10'b0110001000,
    10'b0110000010,
    10'b0101111100,
    10'b0101110110,
    10'b0101110000,
    10'b0101101010,
    10'b0101100100,
    10'b0101011101,
    10'b0101010111,
    10'b0101010000,
    10'b0101001001,
    10'b0101000010,
    10'b0100111011,
    10'b0100110100,
    10'b0100101101,
    10'b0100100110,
    10'b0100011110,
    10'b0100010111,
    10'b0100001111,
    10'b0100001000,
    10'b0100000000,
    10'b0011111000,
    10'b0011110000,
    10'b0011101000,
    10'b0011100000,
    10'b0011011000,
    10'b0011010000,
    10'b0011001000,
    10'b0011000000,
    10'b0010110111,
    10'b0010101111,
    10'b0010100111,
    10'b0010011110,
    10'b0010010110,
    10'b0010001101,
    10'b0010000101,
    10'b0001111100,
    10'b0001110011,
    10'b0001101010,
    10'b0001100010,
    10'b0001011001,
    10'b0001010000,
    10'b0001000111,
    10'b0000111110,
    10'b0000110110,
    10'b0000101101,
    10'b0000100100,
    10'b0000011011,
    10'b0000010010,
    10'b0000001001,
    10'b0000000000,
    10'b1111110111,
    10'b1111101110,
    10'b1111100101,
    10'b1111011100,
    10'b1111010011,
    10'b1111001010,
    10'b1111000010,
    10'b1110111001,
    10'b1110110000,
    10'b1110100111,
    10'b1110011110,
    10'b1110010110,
    10'b1110001101,
    10'b1110000100,
    10'b1101111011,
    10'b1101110011,
    10'b1101101010,
    10'b1101100010,
    10'b1101011001,
    10'b1101010001,
    10'b1101001001,
    10'b1101000000,
    10'b1100111000,
    10'b1100110000,
    10'b1100101000,
    10'b1100100000,
    10'b1100011000,
    10'b1100010000,
    10'b1100001000,
    10'b1100000000,
    10'b1011111000,
    10'b1011110001,
    10'b1011101001,
    10'b1011100010,
    10'b1011011010,
    10'b1011010011,
    10'b1011001100,
    10'b1011000101,
    10'b1010111110,
    10'b1010110111,
    10'b1010110000,
    10'b1010101001,
    10'b1010100011,
    10'b1010011100,
    10'b1010010110,
    10'b1010010000,
    10'b1010001010,
    10'b1010000100,
    10'b1001111110,
    10'b1001111000,
    10'b1001110010,
    10'b1001101101,
    10'b1001100111,
    10'b1001100010,
    10'b1001011101,
    10'b1001011000,
    10'b1001010011,
    10'b1001001110,
    10'b1001001001,
    10'b1001000101,
    10'b1001000000,
    10'b1000111100,
    10'b1000111000,
    10'b1000110100,
    10'b1000110000,
    10'b1000101100,
    10'b1000101001,
    10'b1000100101,
    10'b1000100010,
    10'b1000011111,
    10'b1000011100,
    10'b1000011001,
    10'b1000010110,
    10'b1000010100,
    10'b1000010001,
    10'b1000001111,
    10'b1000001101,
    10'b1000001011,
    10'b1000001001,
    10'b1000001000,
    10'b1000000110,
    10'b1000000101,
    10'b1000000100,
    10'b1000000011,
    10'b1000000010,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000001,
    10'b1000000010,
    10'b1000000011,
    10'b1000000100,
    10'b1000000101,
    10'b1000000110,
    10'b1000001000,
    10'b1000001001,
    10'b1000001011,
    10'b1000001101,
    10'b1000001111,
    10'b1000010001,
    10'b1000010100,
    10'b1000010110,
    10'b1000011001,
    10'b1000011100,
    10'b1000011111,
    10'b1000100010,
    10'b1000100101,
    10'b1000101001,
    10'b1000101100,
    10'b1000110000,
    10'b1000110100,
    10'b1000111000,
    10'b1000111100,
    10'b1001000000,
    10'b1001000101,
    10'b1001001001,
    10'b1001001110,
    10'b1001010011,
    10'b1001011000,
    10'b1001011101,
    10'b1001100010,
    10'b1001100111,
    10'b1001101101,
    10'b1001110010,
    10'b1001111000,
    10'b1001111110,
    10'b1010000100,
    10'b1010001010,
    10'b1010010000,
    10'b1010010110,
    10'b1010011100,
    10'b1010100011,
    10'b1010101001,
    10'b1010110000,
    10'b1010110111,
    10'b1010111110,
    10'b1011000101,
    10'b1011001100,
    10'b1011010011,
    10'b1011011010,
    10'b1011100010,
    10'b1011101001,
    10'b1011110001,
    10'b1011111000,
    10'b1100000000,
    10'b1100001000,
    10'b1100010000,
    10'b1100011000,
    10'b1100100000,
    10'b1100101000,
    10'b1100110000,
    10'b1100111000,
    10'b1101000000,
    10'b1101001001,
    10'b1101010001,
    10'b1101011001,
    10'b1101100010,
    10'b1101101010,
    10'b1101110011,
    10'b1101111011,
    10'b1110000100,
    10'b1110001101,
    10'b1110010110,
    10'b1110011110,
    10'b1110100111,
    10'b1110110000,
    10'b1110111001,
    10'b1111000010,
    10'b1111001010,
    10'b1111010011,
    10'b1111011100,
    10'b1111100101,
    10'b1111101110,
    10'b1111110111
};

reg signed [9:0] dir_x = Dir_x[180]; // * 2 ^ 9
reg signed [9:0] dir_y = Dir_y[180]; // * 2 ^ 9
wire signed [9:0] hor_x;             // * 2 ^ 9
wire signed [9:0] hor_y;             // * 2 ^ 9
assign hor_x = dir_y;
assign hor_y = -dir_x;
/*
R = [[hor_x,    0,   dir_x],
     [hor_y,    0,   dir_y],
     [    0,   -1,       0]]
*/

reg [9:0] tmp[1:0];
reg signed [9:0] ray_dir[2:0];   // * 2 ^ 9
reg signed [9:0] ray_dir_R[1:0][2:0]; // * 2 ^ 8

wire signed [18:0] hor_p_1[5:0];
wire signed [18:0] ver_p_1[5:0];
wire signed [18:0] ground_1;
wire [9:0] hor_p_2[5:0];
wire [9:0] ver_p_2[5:0];
wire [9:0] ground_2;
wire [9:0] hor_p_3[5:0];
wire [9:0] ver_p_3[5:0];
wire [9:0] ground_3;
wire signed [11:0] hor_out_1[5:0][2:0];
wire signed [11:0] ver_out_1[5:0][2:0];
wire signed [11:0] ground_out_1[2:0];
wire signed [9:0] hor_out_2[5:0][2:0];
wire signed [9:0] ver_out_2[5:0][2:0];
wire signed [9:0] ground_out_2[2:0];
wire [5:0] hor_en;
wire [5:0] ver_en;
wire ground_en;

reg outp_en;
reg signed [9:0] outp;
reg rev;
reg [1:0] normal_dir;

wire signed [9:0] dir_to_light[3:0][2:0];

genvar xx;
generate
    for (xx = 0; xx < 6; xx = xx + 1) begin: hor
        intersection #(xx) intersection_x(
            .clk(clk_vga),
            .dir(ray_dir_R[0][0]),
            .ori(center_x),
            .p(hor_p_1[xx])
        );
        get_pos getter_x(
            .clk(clk_vga),
            .p(hor_p_1[xx]),
            .ori_x({1'b0, center_x}),
            .ori_y({1'b0, center_y}),
            .ori_z({1'b0, center_z}),
            .dir_x(ray_dir_R[1][0]),
            .dir_y(ray_dir_R[1][1]),
            .dir_z(ray_dir_R[1][2]),
            .out_x(hor_out_1[xx][0]),
            .out_y(hor_out_1[xx][1]),
            .out_z(hor_out_1[xx][2]),
            .out_p(hor_p_2[xx])
        );
        check_valid #(xx) checker_x(
            .clk(clk_vga),
            .wall(hor_wall[xx]),
            .in_p(hor_p_2[xx]),
            .in_x(hor_out_1[xx][1]),
            .in_y(hor_out_1[xx][2]),
            .in_z(hor_out_1[xx][0]),
            .out_x(hor_out_2[xx][1]),
            .out_y(hor_out_2[xx][2]),
            .out_z(hor_out_2[xx][0]),
            .out_p(hor_p_3[xx]),
            .en(hor_en[xx])
        );
    end
endgenerate

genvar yy;
generate
    for (yy = 0; yy < 6; yy = yy + 1) begin: ver
        intersection #(yy) intersection_y(
            .clk(clk_vga),
            .dir(ray_dir_R[0][1]),
            .ori(center_y),
            .p(ver_p_1[yy])
        );
        get_pos getter_y(
            .clk(clk_vga),
            .p(ver_p_1[yy]),
            .ori_x({1'b0, center_x}),
            .ori_y({1'b0, center_y}),
            .ori_z({1'b0, center_z}),
            .dir_x(ray_dir_R[1][0]),
            .dir_y(ray_dir_R[1][1]),
            .dir_z(ray_dir_R[1][2]),
            .out_x(ver_out_1[yy][0]),
            .out_y(ver_out_1[yy][1]),
            .out_z(ver_out_1[yy][2]),
            .out_p(ver_p_2[yy])
        );
        check_valid #(yy) checker_y(
            .clk(clk_vga),
            .wall(ver_wall[yy]),
            .in_p(ver_p_2[yy]),
            .in_x(ver_out_1[yy][0]),
            .in_y(ver_out_1[yy][2]),
            .in_z(ver_out_1[yy][1]),
            .out_x(ver_out_2[yy][0]),
            .out_y(ver_out_2[yy][2]),
            .out_z(ver_out_2[yy][1]),
            .out_p(ver_p_3[yy]),
            .en(ver_en[yy])
        );
    end
endgenerate

intersection #(0) intersection_z(
    .clk(clk_vga),
    .dir(ray_dir_R[0][2]),
    .ori(center_z),
    .p(ground_1)
);

get_pos getter_z(
    .clk(clk_vga),
    .p(ground_1),
    .ori_x({1'b0, center_x}),
    .ori_y({1'b0, center_y}),
    .ori_z({1'b0, center_z}),
    .dir_x(ray_dir_R[1][0]),
    .dir_y(ray_dir_R[1][1]),
    .dir_z(ray_dir_R[1][2]),
    .out_x(ground_out_1[0]),
    .out_y(ground_out_1[1]),
    .out_z(ground_out_1[2]),
    .out_p(ground_2)
);

check_valid_ground checker_z(
    .clk(clk_vga),
    .in_p(ground_2),
    .in_x(ground_out_1[0]),
    .in_y(ground_out_1[1]),
    .in_z(ground_out_1[2]),
    .out_x(ground_out_2[0]),
    .out_y(ground_out_2[1]),
    .out_z(ground_out_2[2]),
    .out_p(ground_3),
    .en(ground_en)
);

get_min miner(
    .clk(clk_vga),
    .x(x),
    .y(y),
    .p1_en(ground_en),
    .p1(ground_3),
    .p1_x(ground_out_2[0]),
    .p1_y(ground_out_2[1]),
    .p1_z(ground_out_2[2]),
    .p2_en(hor_en[0]),
    .p2(hor_p_3[0]),
    .p2_x(hor_out_2[0][0]),
    .p2_y(hor_out_2[0][1]),
    .p2_z(hor_out_2[0][2]),
    .p3_en(hor_en[1]),
    .p3(hor_p_3[1]),
    .p3_x(hor_out_2[1][0]),
    .p3_y(hor_out_2[1][1]),
    .p3_z(hor_out_2[1][2]),
    .p4_en(hor_en[2]),
    .p4(hor_p_3[2]),
    .p4_x(hor_out_2[2][0]),
    .p4_y(hor_out_2[2][1]),
    .p4_z(hor_out_2[2][2]),
    .p5_en(hor_en[3]),
    .p5(hor_p_3[3]),
    .p5_x(hor_out_2[3][0]),
    .p5_y(hor_out_2[3][1]),
    .p5_z(hor_out_2[3][2]),
    .p6_en(hor_en[4]),
    .p6(hor_p_3[4]),
    .p6_x(hor_out_2[4][0]),
    .p6_y(hor_out_2[4][1]),
    .p6_z(hor_out_2[4][2]),
    .p7_en(hor_en[5]),
    .p7(hor_p_3[5]),
    .p7_x(hor_out_2[5][0]),
    .p7_y(hor_out_2[5][1]),
    .p7_z(hor_out_2[5][2]),
    .p8_en(ver_en[0]),
    .p8(ver_p_3[0]),
    .p8_x(ver_out_2[0][0]),
    .p8_y(ver_out_2[0][1]),
    .p8_z(ver_out_2[0][2]),
    .p9_en(ver_en[1]),
    .p9(ver_p_3[1]),
    .p9_x(ver_out_2[1][0]),
    .p9_y(ver_out_2[1][1]),
    .p9_z(ver_out_2[1][2]),
    .p10_en(ver_en[2]),
    .p10(ver_p_3[2]),
    .p10_x(ver_out_2[2][0]),
    .p10_y(ver_out_2[2][1]),
    .p10_z(ver_out_2[2][2]),
    .p11_en(ver_en[3]),
    .p11(ver_p_3[3]),
    .p11_x(ver_out_2[3][0]),
    .p11_y(ver_out_2[3][1]),
    .p11_z(ver_out_2[3][2]),
    .p12_en(ver_en[4]),
    .p12(ver_p_3[4]),
    .p12_x(ver_out_2[4][0]),
    .p12_y(ver_out_2[4][1]),
    .p12_z(ver_out_2[4][2]),
    .p13_en(ver_en[5]),
    .p13(ver_p_3[5]),
    .p13_x(ver_out_2[5][0]),
    .p13_y(ver_out_2[5][1]),
    .p13_z(ver_out_2[5][2]),
    .outp_en(outp_en),
    .outp(outp),
    .rev(rev),
    .normal_dir(normal_dir), // 0: x 1: y 2: z
    .dir_to_light_0_x(dir_to_light[0][0]),
    .dir_to_light_0_y(dir_to_light[0][1]),
    .dir_to_light_0_z(dir_to_light[0][2]),
    .dir_to_light_1_x(dir_to_light[1][0]),
    .dir_to_light_1_y(dir_to_light[1][1]),
    .dir_to_light_1_z(dir_to_light[1][2]),
    .dir_to_light_2_x(dir_to_light[2][0]),
    .dir_to_light_2_y(dir_to_light[2][1]),
    .dir_to_light_2_z(dir_to_light[2][2]),
    .dir_to_light_3_x(dir_to_light[3][0]),
    .dir_to_light_3_y(dir_to_light[3][1]),
    .dir_to_light_3_z(dir_to_light[3][2])
);

reg [7:0] tmp_comp[2:0];
localparam [0:3][2:0] light_color = {3'b111, 3'b111, 3'b111, 3'b111};
localparam [0:3][23:0] light_color_comp = {{8'd192, 8'd128, 8'd128}, {8'd192, 8'd128, 8'd128}, {8'd192, 8'd128, 8'd128}, {8'd192, 8'd128, 8'd128}};
reg signed [9:0] single_shade[3:0][2:0];
reg signed [9:0] single_shade_comp[3:0][2:0];
reg [7:0] phone[2:0];

reg [7:0] red;
reg [7:0] green;
reg [7:0] blue;
assign wr_data = {{8{1'b0}}, red, green, blue};

reg [31:0] debug/*synthesis noprune*/;
reg [31:0] debug_2/*synthesis noprune*/;
reg [31:0] debug_3/*synthesis noprune*/;
reg [31:0] debug_4/*synthesis noprune*/;

// main states
always @ (posedge clk_vga or posedge reset_btn) begin
    if (reset_btn) begin
        draw_mode <= RIGHT;
        image_cnt <= 8'd90;
        center_angle <= 9'd180;
        {center_x, center_y} <= {10'd32, 10'd32};
        x <= 3'd0;
        y <= 3'd0;
        dir <= D;
        move_en <= 1'b1;
        state <= INIT_CAM;
        enter_state <= COVER_PHASE1;
        grad_rate <= 17'd0;
        wr_en <= 1'b0;
        center_z <= 120;
        // wr_addr <= 19'b0;
        pip_en <= 9'b111111111;
    end
    else begin
        case (state)
            STILL: begin
                if (x == 4 && y == 4) begin
                    grad_rate <= 0;
                    enter_state <= FINAL_PHASE;
                    state <= INIT_CAM;
                end
                else if (!move_en && signal) begin
                    case (move_data)
                        MOVE: begin
                            case (dir)
                                U: begin
                                    if (x > 3'd0 && !maze[x - 1][y]) begin
                                        draw_mode <= move_data;
                                        state <= INIT_CAM;
                                        image_cnt <= 8'd0;
                                    end
                                end
                                L: begin
                                    if (y > 3'd0 && !maze[x][y - 1]) begin
                                        draw_mode <= move_data;
                                        state <= INIT_CAM;
                                        image_cnt <= 8'd0;
                                    end
                                end
                                D: begin
                                    if (x < 3'd4 && !maze[x + 1][y]) begin
                                        draw_mode <= move_data;
                                        state <= INIT_CAM;
                                        image_cnt <= 8'd0;
                                    end
                                end
                                R: begin
                                    if (y < 3'd4 && !maze[x][y + 1]) begin
                                        draw_mode <= move_data;
                                        state <= INIT_CAM;
                                        image_cnt <= 8'd0;
                                    end
                                end
                            endcase
                        end
                        LEFT, RIGHT: begin
                            draw_mode <= move_data;
                            state <= INIT_CAM;
                            image_cnt <= 8'd0;
                        end
                        DARKEN: begin
                            grad_rate <= 17'd0;
                            state <= INIT_CAM;
                            image_cnt <= 8'd0;
                        end
                        UP: begin
                            draw_mode <= move_data;
                            state <= INIT_CAM;
                            image_cnt <= 8'd0;
                        end
                        DOWN: begin
                            draw_mode <= move_data;
                            state <= INIT_CAM;
                            image_cnt <= 8'd0;
                        end
                        default: state <= state;
                    endcase
                    move_en <= 1'b1;
                end
                else if (!signal) begin
                    move_en <= 1'b0;
                end
            end
            INIT_CAM: begin
                //INIT_CAM
                if (!signal) begin
                    move_en <= 1'b0;
                end
                px[0] <= 10'd0;
                px[1] <= 10'd0;
                px[2] <= 10'd0;
                px[3] <= 10'd0;
                px[4] <= 10'd0;
                px[5] <= 10'd0;
                px[6] <= 10'd0;
                px[7] <= 10'd0;
                px[8] <= 10'd0;
                py[0] <= height - 1;
                py[1] <= height - 1;
                py[2] <= height - 1;
                py[3] <= height - 1;
                py[4] <= height - 1;
                py[5] <= height - 1;
                py[6] <= height - 1;
                py[7] <= height - 1;
                py[8] <= height - 1;
                pip_en <= 9'b111111111;
                wr_addr <= 19'b0;
                wr_en <= 1'b0;
                if (enter_state == COVER_PHASE1) begin
                    if (grad_rate < 256) begin
                        grad_rate <= grad_rate + 1;
                    end
                    else begin
                        enter_state <= COVER_PHASE2;
                    end

                    state <= DRAW;
                end
                else if (enter_state == COVER_PHASE2) begin
                    if (grad_rate > 0) begin
                        grad_rate <= grad_rate - 1;
                    end
                    else begin
                        enter_state <= ENTER_PHASE1;
                    end

                    state <= DRAW;
                end
                else if (enter_state == FINAL_PHASE) begin
                    if (grad_rate < 256) begin
                        grad_rate <= grad_rate + 1;
                    end

                    state <= DRAW;
                end
                else if (enter_state == ENTER_PHASE1) begin
                    if (center_y < 287) begin
                        center_y <= center_y + 1;
                        grad_rate <= grad_rate + 1;
                    end
                    else begin
                        center_y <= center_y + 1;
                        grad_rate <= 0;
                        center_angle <= 270;
                        enter_state <= ENTER_PHASE2;
                    end

                    state <= DRAW;
                end
                else if (enter_state == ENTER_PHASE2) begin
                    if (center_x < 287) begin
                        center_x <= center_x + 1;
                        grad_rate <= grad_rate + 1;
                    end
                    else begin
                        center_x <= center_x + 1;
                        grad_rate <= 0;
                        center_x <= 32;
                        center_y <= 32;
                        center_angle <= 180;
                        enter_state <= ENTER_PHASE3;
                    end

                    state <= DRAW;
                end
                else if (enter_state == ENTER_PHASE3) begin
                    if (grad_rate < 258) begin
                        grad_rate <= grad_rate + 4;
                        state <= DRAW;
                    end
                    else if (center_z > 48) begin
                        grad_rate <= 258;
                        center_z <= center_z - 1;
                        state <= DRAW;
                    end
                    else begin
                        enter_state <= NONE;
                        state <= STILL;
                    end
                end
                else if (grad_rate < 17'd256) begin
                    grad_rate <= grad_rate + 2;
                    state <= DRAW;
                end
                else if (grad_rate == 17'd256) begin
                    grad_rate <= grad_rate + 2;
                    state <= STILL;
                end
                else if (draw_mode == UP) begin
                    if (center_z != 288 && image_cnt < 8'd24) begin
                        center_z <= center_z + 1;
                        image_cnt <= image_cnt + 1;
                        state <= DRAW;
                    end
                    else begin
                        image_cnt <= 8'd0;
                        state <= STILL;
                    end
                end
                else if (draw_mode == DOWN) begin
                    if (center_z != 24 && image_cnt < 8'd24) begin
                        center_z <= center_z - 1;
                        image_cnt <= image_cnt + 1;
                        state <= DRAW;
                    end
                    else begin
                        image_cnt <= 8'd0;
                        state <= STILL;
                    end
                end
                else if ((image_cnt == 8'd90 && (draw_mode == LEFT || draw_mode == RIGHT)) || (image_cnt == unit_size && draw_mode == MOVE)) begin
                    image_cnt <= 8'd0;
                    state <= STILL;
                    case (draw_mode)
                        MOVE:
                            case (dir)
                                U: begin
                                    if (x > 3'd0 && !maze[x - 1][y])
                                        x <= x - 1;
                                end
                                L: begin
                                    if (y > 3'd0 && !maze[x][y - 1])
                                        y <= y - 1;
                                end
                                D: begin
                                    if (x < 3'd4 && !maze[x + 1][y])
                                        x <= x + 1;
                                end
                                R: begin
                                    if (y < 3'd4 && !maze[x][y + 1])
                                        y <= y + 1;
                                end
                            endcase
                        LEFT, RIGHT:
                            case (dir)
                                U: begin
                                    if (draw_mode == LEFT)
                                        dir <= L;
                                    else
                                        dir <= R;
                                end
                                L: begin
                                    if (draw_mode == LEFT)
                                        dir <= D;
                                    else
                                        dir <= U;
                                end
                                D: begin
                                    if (draw_mode == LEFT)
                                        dir <= R;
                                    else
                                        dir <= L;
                                end
                                R: begin
                                    if (draw_mode == LEFT)
                                        dir <= U;
                                    else
                                        dir <= D;
                                end
                                endcase
                    endcase
                end
                else begin
                    image_cnt <= image_cnt + 1'b1;
                    state <= DRAW;
                    case (draw_mode)
                        MOVE:
                            case (dir)
                                U: begin
                                    center_x <= center_x - 1;
                                    center_y <= center_y;
                                end
                                L: begin
                                    center_x <= center_x;
                                    center_y <= center_y - 1;
                                end
                                D: begin
                                    center_x <= center_x + 1;
                                    center_y <= center_y;
                                end
                                R: begin
                                    center_x <= center_x;
                                    center_y <= center_y + 1;
                                end
                            endcase
                        LEFT: begin
                            if (center_angle == 9'd0)
                                center_angle <= 9'd359;
                            else
                                center_angle <= center_angle - 1;
                        end
                        RIGHT: begin
                            if (center_angle == 9'd359)
                                center_angle <= 9'd0;
                            else
                                center_angle <= center_angle + 1;
                        end
                    endcase
                end
            end
            DRAW: begin
                dir_x <= Dir_x[center_angle];
                dir_y <= Dir_y[center_angle];
                // 流水线
                if (!signal) begin
                    move_en <= 1'b0;
                end
                px[1] <= px[0];
                px[2] <= px[1];
                px[3] <= px[2];
                px[4] <= px[3];
                px[5] <= px[4];
                px[6] <= px[5];
                px[7] <= px[6];
                px[8] <= px[7];

                py[1] <= py[0];
                py[2] <= py[1];
                py[3] <= py[2];
                py[4] <= py[3];
                py[5] <= py[4];
                py[6] <= py[5];
                py[7] <= py[6];
                py[8] <= py[7];

                pip_en[1] <= pip_en[0];
                pip_en[2] <= pip_en[1];
                pip_en[3] <= pip_en[2];
                pip_en[4] <= pip_en[3];
                pip_en[5] <= pip_en[4];
                pip_en[6] <= pip_en[5];
                pip_en[7] <= pip_en[6];
                pip_en[8] <= pip_en[7];

                ray_dir_R[1] <= ray_dir_R[0];

                // GEN_RAY 1
                if (pip_en[0] == 1'b1) begin // 激活
                    if (px[0] == width) begin
                        pip_en[0] <= 1'b1;
                        px[0] <= width;
                        py[0] <= height;
                    end
                    else begin
                        pip_en[0] <= 1'b0;
                        px[0] <= 10'd0;
                        py[0] <= height - 1;
                        ray_dir[0] <= -400;
                        ray_dir[1] <= -300;
                        ray_dir[2] <= 511;
                    end
                end
                else begin
                    if (px[0] == width - 1 && py[0] == 0) begin
                        pip_en[0] <= 1'b1;
                        px[0] <= width;
                        py[0] <= height;
                    end
                    else if (px[0] == width - 1) begin
                        pip_en[0] <= 1'b0;
                        px[0] <= 10'd0;
                        py[0] <= py[0] - 1;
                        ray_dir[0] <= -400;
                        ray_dir[1] <= 301 - py[0];
                        ray_dir[2] <= 511;
                    end
                    else begin
                        pip_en[0] <= 1'b0;
                        px[0] <= px[0] + 1;
                        py[0] <= py[0];
                        ray_dir[0] <= px[0] - 399;
                        ray_dir[1] <= 300 - py[0];
                        ray_dir[2] <= 511;
                    end
                end

                // GEN_RAY 2
                if (pip_en[0] == 1'b0) begin
                    // do GEN_RAY
                    {ray_dir_R[0][0], tmp[0]} <= ray_dir[0] * hor_x
                                               + ray_dir[2] * dir_x;
                    {ray_dir_R[0][1], tmp[1]} <= ray_dir[0] * hor_y
                                               + ray_dir[2] * dir_y;
                    ray_dir_R[0][2] <= -(ray_dir[1] / 2);
                end
                else begin
                    // stay
                end
                
                // if (px[2] == 600 && py[2] == 150 && center_angle == 180 && center_x == 32 && center_y == 32) begin
                //     debug[18:0] <= hor_p_1[0];
                //     debug_2[9:0] <= ray_dir_R[1][0];
                //     debug_3[9:0] <= ray_dir_R[1][1];
                // end

                if (px[3] == 600 && py[3] == 150 && center_angle == 180 && center_x == 32 && center_y == 32) begin
                    debug[11:0] <= ver_out_1[0][0];
                    debug_2[11:0] <= ver_out_1[0][1];
                    debug_3[11:0] <= ver_out_1[0][2];
                end

                // INTERSECT 1
                if (pip_en[1] == 1'b0) begin
                    // do intersect
                end
                else begin
                    // stay
                end

                // INTERSECT 2
                if (pip_en[2] == 1'b0) begin
                    // do intersect
                end
                else begin
                    // stay
                end

                // INTERSECT 3
                if (pip_en[3] == 1'b0) begin
                    // do intersect
                end
                else begin
                    // stay
                end

                // INTERSECT 4
                if (pip_en[4] == 1'b0) begin
                    // do intersect
                end
                else begin
                    // stay
                end

                // PHONG 1
                if (pip_en[5] == 1'b0) begin
                    // do phong
                    integer i;
                    integer j;
                    if (rev) begin
                        for (i = 0; i < 4; i = i + 1) begin
                            for (j = 0; j < 3; j = j + 1)
                                single_shade[i][j] <= light_color[i][j] ? -dir_to_light[i][normal_dir] : 0;
                            {single_shade_comp[i][0], tmp_comp[0]} <= (-dir_to_light[i][normal_dir] * light_color_comp[i][23:16]);
                            {single_shade_comp[i][1], tmp_comp[1]} <= (-dir_to_light[i][normal_dir] * light_color_comp[i][15:8]);
                            {single_shade_comp[i][2], tmp_comp[2]} <= (-dir_to_light[i][normal_dir] * light_color_comp[i][7:0]);
                        end
                    end
                    else begin
                        for (i = 0; i < 4; i = i + 1) begin
                            for (j = 0; j < 3; j = j + 1)
                                single_shade[i][j] <= light_color[i][j] ? dir_to_light[i][normal_dir] : 0;
                            {single_shade_comp[i][0], tmp_comp[0]} <= (dir_to_light[i][normal_dir] * light_color_comp[i][23:16]);
                            {single_shade_comp[i][1], tmp_comp[1]} <= (dir_to_light[i][normal_dir] * light_color_comp[i][15:8]);
                            {single_shade_comp[i][2], tmp_comp[2]} <= (dir_to_light[i][normal_dir] * light_color_comp[i][7:0]);
                        end
                    end
                end
                else begin
                    // stay
                end

                // PHONG 2
                if (pip_en[6] == 1'b0) begin
                    // do phong
                    if (enter_state == COVER_PHASE1 || enter_state == COVER_PHASE2 || enter_state == FINAL_PHASE) begin
                        if (px[6] < 200 || px[6] > 599 || py[6] < 150 || py[6] > 449) begin
                            phone[0] <= (grad_rate * 16'd255) >> 8;
                            phone[1] <= (grad_rate * 16'd255) >> 8;
                            phone[2] <= (grad_rate * 16'd255) >> 8;
                        end
                        else begin
                            if (enter_state == COVER_PHASE1 || enter_state == COVER_PHASE2) begin
                                phone[0] <= (grad_rate * start_img[15'b0 + ((px[6] - 200) >> 2) + (((449 - py[6]) >> 2) * 100)][23:16]) >> 8;
                                phone[1] <= (grad_rate * start_img[15'b0 + ((px[6] - 200) >> 2) + (((449 - py[6]) >> 2) * 100)][15:8]) >> 8;
                                phone[2] <= (grad_rate * start_img[15'b0 + ((px[6] - 200) >> 2) + (((449 - py[6]) >> 2) * 100)][7:0]) >> 8;
                            end
                            else begin
                                phone[0] <= (grad_rate * end_img[15'b0 + ((px[6] - 200) >> 2) + (((449 - py[6]) >> 2) * 100)][23:16]) >> 8;
                                phone[1] <= (grad_rate * end_img[15'b0 + ((px[6] - 200) >> 2) + (((449 - py[6]) >> 2) * 100)][15:8]) >> 8;
                                phone[2] <= (grad_rate * end_img[15'b0 + ((px[6] - 200) >> 2) + (((449 - py[6]) >> 2) * 100)][7:0]) >> 8;
                            end
                        end
                    end
                    else if (~outp_en) begin
                        if (grad_rate < 17'd258) begin
                            phone[0] <= (grad_rate * 16'd87) >> 8;
                            phone[1] <= (grad_rate * 16'd250) >> 8;
                            phone[2] <= (grad_rate * 16'd255) >> 8;
                        end
                        else begin
                            phone[0] <= 8'd87;
                            phone[1] <= 8'd250;
                            phone[2] <= 8'd255;
                        end
                        
                    end
                    else begin
                        integer i;
                        for (i = 0; i < 3; i = i + 1)
                            // phone[i] <= ((single_shade[0][i][9] ? 0 : single_shade[0][i])
                            //            + (single_shade[1][i][9] ? 0 : single_shade[1][i])
                            //            + (single_shade[2][i][9] ? 0 : single_shade[2][i])
                            //            + (single_shade[3][i][9] ? 0 : single_shade[3][i])) >> 3;
                            if (grad_rate < 17'd258) begin
                                phone[i] <= (grad_rate * (((single_shade_comp[0][i][9] ? 0 : single_shade_comp[0][i])
                                       + (single_shade_comp[1][i][9] ? 0 : single_shade_comp[1][i])
                                       + (single_shade_comp[2][i][9] ? 0 : single_shade_comp[2][i])
                                       + (single_shade_comp[3][i][9] ? 0 : single_shade_comp[3][i])) >> 3)) >> 8;
                            end
                            else begin
                                phone[i] <= ((single_shade_comp[0][i][9] ? 0 : single_shade_comp[0][i])
                                       + (single_shade_comp[1][i][9] ? 0 : single_shade_comp[1][i])
                                       + (single_shade_comp[2][i][9] ? 0 : single_shade_comp[2][i])
                                       + (single_shade_comp[3][i][9] ? 0 : single_shade_comp[3][i])) >> 3;
                            end

                    end
                end
                else begin
                    // stay
                end

                // SET_PIXEL
                if (pip_en[7] == 1'b0) begin
                    // do set_pixel
                    wr_en <= 1'b1;
                    red <= phone[0];
                    green <= phone[1];
                    blue <= phone[2];
                    // red <= px[6];
                    // green <= 100;
                    // blue <= 100;
                end
                else begin
                    // stay
                    wr_en <= 1'b0;
                end

                // back to init_cam
                if (pip_en[8] == 1'b0) begin
                    state <= DRAW;
                end
                else if (px[8] == width) begin
                    state <= INIT_CAM;
                end
                else begin
                    state <= DRAW;
                end

                if (wr_en) begin
                    if (wr_addr == 19'd479999) begin
                        wr_addr <= 19'd0;
                        offset_reg <= offset_reg + 1;
                        // rd_addr_offset <= !rd_addr_offset;
                        // wr_addr_offset <= !wr_addr_offset;
                    end
                    else begin
                        wr_addr <= wr_addr + 1'b1;
                    end
                end
            end
            default:;
        endcase        
    end
    
end

assign video_clk = clk_ps2;
render image_render(
    .clk(clk_100m),
    .clk_vga(clk_vga),
    .clk_50m(clk_ps2),

    .ram_data(base_ram_data),
    .ram_addr(base_ram_addr),
    .ram_ce_n(base_ram_ce_n),
    .ram_oe_n(base_ram_oe_n),
    .ram_we_n(base_ram_we_n),

    .rd_addr_offset(rd_addr_offset),
    .wr_addr_offset(wr_addr_offset),
    .sram_wr_en(wr_en),
    .sram_wr_addr(wr_addr),
    .sram_wr_data(wr_data),

    .vga_hsync(video_hsync),
    .vga_vsync(video_vsync),

    .vga_red(video_red), 
    .vga_green(video_green),
    .vga_blue(video_blue),

    .vga_data_en(video_de)
);
/* =========== Demo code end =========== */

endmodule
